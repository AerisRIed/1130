/*
 * This empty include file is generated and `included in the compile flow.
 * This allows you to create your own file (of the same name) in your own
 * directory and `include your dut_usb4_tc_noc_env_pkg extensions.
 *
 * Your own files can be included in the compile flow by:
 * 1. create <my extensions dir>/env_pkg/dut_usb4_tc_noc_env_pkg_usr.sv
 *    > `include your own TB package extensions files
 * 2. include <my extensions dir>/env_pkg in the compile flow
 *    > stg -sim ... -irunopts "-incdir <my extensions dir>/env_pkg" ...
 *    or 
 *    > irun ... -incdir <my extensions dir>/env_pkg ...
 *
 */
