`ifndef TEST_MAIN__SV
`define TEST_MAIN__SV

`endif