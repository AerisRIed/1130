`include"cdn_message_bus_test.sv"
