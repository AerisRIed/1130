class passive_slave_usb4_tc_noc_apb_mstr_config extends cdnApbUvmConfig;

   `uvm_object_utils(passive_slave_usb4_tc_noc_apb_mstr_config)

   function new(string name = "passive_slave_usb4_tc_noc_apb_mstr_config");
      super.new(name);
   endfunction : new

   virtual function void setFieldsValues();
      set_use_apb_amba4_extension(1);
      set_number_of_slaves(1);
      set_DeviceType(CDN_APB_CFG_SLAVE);
      set_idle_mode_optimization(CDN_APB_CFG_IDLE_MODE_OPTIMIZATION_OPTIMIZED_CB);
      set_is_active(UVM_PASSIVE);
      set_use_apb_ver_d_extension(1);
      set_use_memory(0);

   endfunction: setFieldsValues

endclass : passive_slave_usb4_tc_noc_apb_mstr_config
