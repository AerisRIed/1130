// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc (
  input  wire            tap2apb_pclk,
  input  wire            noc_clk,
  input  wire            rst_n,
  // apb_mstr
  input  wire     [31:0] apb_mstr_paddr,                                        // Address
  input  wire            apb_mstr_psel,                                         // Select
  input  wire            apb_mstr_penable,                                      // Enable
  input  wire            apb_mstr_pwrite,                                       // Write not read
  input  wire     [31:0] apb_mstr_pwdata,                                       // Write data
  input  wire      [3:0] apb_mstr_pstrb,                                        // Write strobes
  output logic           apb_mstr_pready,                                       // Ready
  output logic    [31:0] apb_mstr_prdata,                                       // Read data
  output logic           apb_mstr_pslverr,                                      // Slave error
  // cdb
  input  wire     [31:0] cdb_paddr,                                             // Address
  input  wire            cdb_psel,                                              // Select
  input  wire            cdb_penable,                                           // Enable
  input  wire            cdb_pwrite,                                            // Write not read
  input  wire     [31:0] cdb_pwdata,                                            // Write data
  input  wire      [3:0] cdb_pstrb,                                             // Write strobes
  output logic           cdb_pready,                                            // Ready
  output logic    [31:0] cdb_prdata,                                            // Read data
  output logic           cdb_pslverr,                                           // Slave error
  // cmn_cdb
  output logic     [8:0] cmn_cdb_paddr,                                         // Address
  output logic           cmn_cdb_psel,                                          // Select
  output logic           cmn_cdb_penable,                                       // Enable
  output logic           cmn_cdb_pwrite,                                        // Write not read
  output logic    [31:0] cmn_cdb_pwdata,                                        // Write data
  output logic     [3:0] cmn_cdb_pstrb,                                         // Write strobes
  input  wire            cmn_cdb_pready,                                        // Ready
  input  wire     [31:0] cmn_cdb_prdata,                                        // Read data
  // tc_reg
  output logic    [15:0] tc_reg_paddr,                                          // Address
  output logic           tc_reg_psel,                                           // Select
  output logic           tc_reg_penable,                                        // Enable
  output logic           tc_reg_pwrite,                                         // Write not read
  output logic    [31:0] tc_reg_pwdata,                                         // Write data
  output logic     [3:0] tc_reg_pstrb,                                          // Write strobes
  input  wire            tc_reg_pready,                                         // Ready
  input  wire     [31:0] tc_reg_prdata,                                         // Read data
  // usb_sub_sys
  output logic    [15:0] usb_sub_sys_paddr,                                     // Address
  output logic           usb_sub_sys_psel,                                      // Select
  output logic           usb_sub_sys_penable,                                   // Enable
  output logic           usb_sub_sys_pwrite,                                    // Write not read
  output logic    [31:0] usb_sub_sys_pwdata,                                    // Write data
  output logic     [3:0] usb_sub_sys_pstrb,                                     // Write strobes
  input  wire            usb_sub_sys_pready,                                    // Ready
  input  wire     [31:0] usb_sub_sys_prdata,                                    // Read data
  // pam3_sub_sys
  output logic    [15:0] pam3_sub_sys_paddr,                                    // Address
  output logic           pam3_sub_sys_psel,                                     // Select
  output logic           pam3_sub_sys_penable,                                  // Enable
  output logic           pam3_sub_sys_pwrite,                                   // Write not read
  output logic    [31:0] pam3_sub_sys_pwdata,                                   // Write data
  output logic     [3:0] pam3_sub_sys_pstrb,                                    // Write strobes
  input  wire            pam3_sub_sys_pready,                                   // Ready
  input  wire     [31:0] pam3_sub_sys_prdata,                                   // Read data
  // apb_tgt
  output logic    [17:0] apb_tgt_paddr,                                         // Address
  output logic           apb_tgt_psel,                                          // Select
  output logic           apb_tgt_penable,                                       // Enable
  output logic           apb_tgt_pwrite,                                        // Write not read
  output logic    [31:0] apb_tgt_pwdata,                                        // Write data
  output logic     [3:0] apb_tgt_pstrb,                                         // Write strobes
  input  wire            apb_tgt_pready,                                        // Ready
  input  wire     [31:0] apb_tgt_prdata,                                        // Read data
  input  wire            apb_tgt_pslverr,                                       // Slave error
  // xcvr_ln_0
  output logic     [9:0] xcvr_ln_0_paddr,                                       // Address
  output logic           xcvr_ln_0_psel,                                        // Select
  output logic           xcvr_ln_0_penable,                                     // Enable
  output logic           xcvr_ln_0_pwrite,                                      // Write not read
  output logic    [31:0] xcvr_ln_0_pwdata,                                      // Write data
  output logic     [3:0] xcvr_ln_0_pstrb,                                       // Write strobes
  input  wire            xcvr_ln_0_pready,                                      // Ready
  input  wire     [31:0] xcvr_ln_0_prdata                                       // Read data
);

logic           apb_mstr_f0_activity;                                           // Upcoming activity indicator
logic           apb_mstr_f0_req;                                                // Flit transfer request
logic           apb_mstr_f0_sop;                                                // Start of packet indicator
logic           apb_mstr_f0_eop;                                                // End of packet indicator
logic    [35:0] apb_mstr_f0_flitdata;                                           // Flit data
logic           apb_mstr_f0_ready;                                              // Flit transfer ready
logic           apb_mstr_f1_activity;                                           // Upcoming activity indicator
logic           apb_mstr_f1_req;                                                // Flit transfer request
logic           apb_mstr_f1_sop;                                                // Start of packet indicator
logic           apb_mstr_f1_eop;                                                // End of packet indicator
logic    [59:0] apb_mstr_f1_flitdata;                                           // Flit data
logic           apb_mstr_f1_ready;                                              // Flit transfer ready
logic           tap2apb_f0_activity;                                            // Upcoming activity indicator
logic           tap2apb_f0_req;                                                 // Flit transfer request
logic           tap2apb_f0_sop;                                                 // Start of packet indicator
logic           tap2apb_f0_eop;                                                 // End of packet indicator
logic    [35:0] tap2apb_f0_flitdata;                                            // Flit data
logic           tap2apb_f0_ready;                                               // Flit transfer ready
logic           tap2apb_f1_activity;                                            // Upcoming activity indicator
logic           tap2apb_f1_req;                                                 // Flit transfer request
logic           tap2apb_f1_sop;                                                 // Start of packet indicator
logic           tap2apb_f1_eop;                                                 // End of packet indicator
logic    [59:0] tap2apb_f1_flitdata;                                            // Flit data
logic           tap2apb_f1_ready;                                               // Flit transfer ready
logic           pam3_cmn_TEA_r0_activity;                                       // Upcoming activity indicator
logic           pam3_cmn_TEA_r0_req;                                            // Flit transfer request
logic           pam3_cmn_TEA_r0_sop;                                            // Start of packet indicator
logic           pam3_cmn_TEA_r0_eop;                                            // End of packet indicator
logic    [33:0] pam3_cmn_TEA_r0_flitdata;                                       // Flit data
logic           pam3_cmn_TEA_r0_ready;                                          // Flit transfer ready
logic           pam3_cmn_TEA_r1_activity;                                       // Upcoming activity indicator
logic           pam3_cmn_TEA_r1_req;                                            // Flit transfer request
logic           pam3_cmn_TEA_r1_sop;                                            // Start of packet indicator
logic           pam3_cmn_TEA_r1_eop;                                            // End of packet indicator
logic    [23:0] pam3_cmn_TEA_r1_flitdata;                                       // Flit data
logic           pam3_cmn_TEA_r1_ready;                                          // Flit transfer ready
logic           tc_reg_TEA_r0_activity;                                         // Upcoming activity indicator
logic           tc_reg_TEA_r0_req;                                              // Flit transfer request
logic           tc_reg_TEA_r0_sop;                                              // Start of packet indicator
logic           tc_reg_TEA_r0_eop;                                              // End of packet indicator
logic    [33:0] tc_reg_TEA_r0_flitdata;                                         // Flit data
logic           tc_reg_TEA_r0_ready;                                            // Flit transfer ready
logic           tc_reg_TEA_r1_activity;                                         // Upcoming activity indicator
logic           tc_reg_TEA_r1_req;                                              // Flit transfer request
logic           tc_reg_TEA_r1_sop;                                              // Start of packet indicator
logic           tc_reg_TEA_r1_eop;                                              // End of packet indicator
logic    [23:0] tc_reg_TEA_r1_flitdata;                                         // Flit data
logic           tc_reg_TEA_r1_ready;                                            // Flit transfer ready
logic           usb_sub_sys_TEA_r0_activity;                                    // Upcoming activity indicator
logic           usb_sub_sys_TEA_r0_req;                                         // Flit transfer request
logic           usb_sub_sys_TEA_r0_sop;                                         // Start of packet indicator
logic           usb_sub_sys_TEA_r0_eop;                                         // End of packet indicator
logic    [33:0] usb_sub_sys_TEA_r0_flitdata;                                    // Flit data
logic           usb_sub_sys_TEA_r0_ready;                                       // Flit transfer ready
logic           usb_sub_sys_TEA_r1_activity;                                    // Upcoming activity indicator
logic           usb_sub_sys_TEA_r1_req;                                         // Flit transfer request
logic           usb_sub_sys_TEA_r1_sop;                                         // Start of packet indicator
logic           usb_sub_sys_TEA_r1_eop;                                         // End of packet indicator
logic    [23:0] usb_sub_sys_TEA_r1_flitdata;                                    // Flit data
logic           usb_sub_sys_TEA_r1_ready;                                       // Flit transfer ready
logic           pam3_sub_sys_TEA_r0_activity;                                   // Upcoming activity indicator
logic           pam3_sub_sys_TEA_r0_req;                                        // Flit transfer request
logic           pam3_sub_sys_TEA_r0_sop;                                        // Start of packet indicator
logic           pam3_sub_sys_TEA_r0_eop;                                        // End of packet indicator
logic    [33:0] pam3_sub_sys_TEA_r0_flitdata;                                   // Flit data
logic           pam3_sub_sys_TEA_r0_ready;                                      // Flit transfer ready
logic           pam3_sub_sys_TEA_r1_activity;                                   // Upcoming activity indicator
logic           pam3_sub_sys_TEA_r1_req;                                        // Flit transfer request
logic           pam3_sub_sys_TEA_r1_sop;                                        // Start of packet indicator
logic           pam3_sub_sys_TEA_r1_eop;                                        // End of packet indicator
logic    [23:0] pam3_sub_sys_TEA_r1_flitdata;                                   // Flit data
logic           pam3_sub_sys_TEA_r1_ready;                                      // Flit transfer ready
logic           usb4_phy_TEA_r0_activity;                                       // Upcoming activity indicator
logic           usb4_phy_TEA_r0_req;                                            // Flit transfer request
logic           usb4_phy_TEA_r0_sop;                                            // Start of packet indicator
logic           usb4_phy_TEA_r0_eop;                                            // End of packet indicator
logic    [33:0] usb4_phy_TEA_r0_flitdata;                                       // Flit data
logic           usb4_phy_TEA_r0_ready;                                          // Flit transfer ready
logic           usb4_phy_TEA_r1_activity;                                       // Upcoming activity indicator
logic           usb4_phy_TEA_r1_req;                                            // Flit transfer request
logic           usb4_phy_TEA_r1_sop;                                            // Start of packet indicator
logic           usb4_phy_TEA_r1_eop;                                            // End of packet indicator
logic    [23:0] usb4_phy_TEA_r1_flitdata;                                       // Flit data
logic           usb4_phy_TEA_r1_ready;                                          // Flit transfer ready
logic           pam3_xcvr_TEA_r0_activity;                                      // Upcoming activity indicator
logic           pam3_xcvr_TEA_r0_req;                                           // Flit transfer request
logic           pam3_xcvr_TEA_r0_sop;                                           // Start of packet indicator
logic           pam3_xcvr_TEA_r0_eop;                                           // End of packet indicator
logic    [33:0] pam3_xcvr_TEA_r0_flitdata;                                      // Flit data
logic           pam3_xcvr_TEA_r0_ready;                                         // Flit transfer ready
logic           pam3_xcvr_TEA_r1_activity;                                      // Upcoming activity indicator
logic           pam3_xcvr_TEA_r1_req;                                           // Flit transfer request
logic           pam3_xcvr_TEA_r1_sop;                                           // Start of packet indicator
logic           pam3_xcvr_TEA_r1_eop;                                           // End of packet indicator
logic    [23:0] pam3_xcvr_TEA_r1_flitdata;                                      // Flit data
logic           pam3_xcvr_TEA_r1_ready;                                         // Flit transfer ready
logic           tap2apb_r0_activity;                                            // Upcoming activity indicator
logic           tap2apb_r0_req;                                                 // Flit transfer request
logic           tap2apb_r0_sop;                                                 // Start of packet indicator
logic           tap2apb_r0_eop;                                                 // End of packet indicator
logic    [33:0] tap2apb_r0_flitdata;                                            // Flit data
logic           tap2apb_r0_ready;                                               // Flit transfer ready
logic           tap2apb_r1_activity;                                            // Upcoming activity indicator
logic           tap2apb_r1_req;                                                 // Flit transfer request
logic           tap2apb_r1_sop;                                                 // Start of packet indicator
logic           tap2apb_r1_eop;                                                 // End of packet indicator
logic    [23:0] tap2apb_r1_flitdata;                                            // Flit data
logic           tap2apb_r1_ready;                                               // Flit transfer ready
logic           RTR_INI0_f0_activity;                                           // Upcoming activity indicator
logic           RTR_INI0_f0_req;                                                // Flit transfer request
logic           RTR_INI0_f0_sop;                                                // Start of packet indicator
logic           RTR_INI0_f0_eop;                                                // End of packet indicator
logic    [35:0] RTR_INI0_f0_flitdata;                                           // Flit data
logic           RTR_INI0_f0_ready;                                              // Flit transfer ready
logic           RTR_INI0_f1_activity;                                           // Upcoming activity indicator
logic           RTR_INI0_f1_req;                                                // Flit transfer request
logic           RTR_INI0_f1_sop;                                                // Start of packet indicator
logic           RTR_INI0_f1_eop;                                                // End of packet indicator
logic    [59:0] RTR_INI0_f1_flitdata;                                           // Flit data
logic           RTR_INI0_f1_ready;                                              // Flit transfer ready
logic           apb_mstr_r0_activity;                                           // Upcoming activity indicator
logic           apb_mstr_r0_req;                                                // Flit transfer request
logic           apb_mstr_r0_sop;                                                // Start of packet indicator
logic           apb_mstr_r0_eop;                                                // End of packet indicator
logic    [33:0] apb_mstr_r0_flitdata;                                           // Flit data
logic           apb_mstr_r0_ready;                                              // Flit transfer ready
logic           apb_mstr_r1_activity;                                           // Upcoming activity indicator
logic           apb_mstr_r1_req;                                                // Flit transfer request
logic           apb_mstr_r1_sop;                                                // Start of packet indicator
logic           apb_mstr_r1_eop;                                                // End of packet indicator
logic    [23:0] apb_mstr_r1_flitdata;                                           // Flit data
logic           apb_mstr_r1_ready;                                              // Flit transfer ready
logic           RTR_INI0_r0_activity;                                           // Upcoming activity indicator
logic           RTR_INI0_r0_req;                                                // Flit transfer request
logic           RTR_INI0_r0_sop;                                                // Start of packet indicator
logic           RTR_INI0_r0_eop;                                                // End of packet indicator
logic    [33:0] RTR_INI0_r0_flitdata;                                           // Flit data
logic           RTR_INI0_r0_ready;                                              // Flit transfer ready
logic           RTR_INI0_r1_activity;                                           // Upcoming activity indicator
logic           RTR_INI0_r1_req;                                                // Flit transfer request
logic           RTR_INI0_r1_sop;                                                // Start of packet indicator
logic           RTR_INI0_r1_eop;                                                // End of packet indicator
logic    [23:0] RTR_INI0_r1_flitdata;                                           // Flit data
logic           RTR_INI0_r1_ready;                                              // Flit transfer ready
logic           pam3_cmn_TEA_f0_activity;                                       // Upcoming activity indicator
logic           pam3_cmn_TEA_f0_req;                                            // Flit transfer request
logic           pam3_cmn_TEA_f0_sop;                                            // Start of packet indicator
logic           pam3_cmn_TEA_f0_eop;                                            // End of packet indicator
logic    [35:0] pam3_cmn_TEA_f0_flitdata;                                       // Flit data
logic           pam3_cmn_TEA_f0_ready;                                          // Flit transfer ready
logic           pam3_cmn_TEA_f1_activity;                                       // Upcoming activity indicator
logic           pam3_cmn_TEA_f1_req;                                            // Flit transfer request
logic           pam3_cmn_TEA_f1_sop;                                            // Start of packet indicator
logic           pam3_cmn_TEA_f1_eop;                                            // End of packet indicator
logic    [59:0] pam3_cmn_TEA_f1_flitdata;                                       // Flit data
logic           pam3_cmn_TEA_f1_ready;                                          // Flit transfer ready
logic           tc_reg_TEA_f0_activity;                                         // Upcoming activity indicator
logic           tc_reg_TEA_f0_req;                                              // Flit transfer request
logic           tc_reg_TEA_f0_sop;                                              // Start of packet indicator
logic           tc_reg_TEA_f0_eop;                                              // End of packet indicator
logic    [35:0] tc_reg_TEA_f0_flitdata;                                         // Flit data
logic           tc_reg_TEA_f0_ready;                                            // Flit transfer ready
logic           tc_reg_TEA_f1_activity;                                         // Upcoming activity indicator
logic           tc_reg_TEA_f1_req;                                              // Flit transfer request
logic           tc_reg_TEA_f1_sop;                                              // Start of packet indicator
logic           tc_reg_TEA_f1_eop;                                              // End of packet indicator
logic    [59:0] tc_reg_TEA_f1_flitdata;                                         // Flit data
logic           tc_reg_TEA_f1_ready;                                            // Flit transfer ready
logic           usb_sub_sys_TEA_f0_activity;                                    // Upcoming activity indicator
logic           usb_sub_sys_TEA_f0_req;                                         // Flit transfer request
logic           usb_sub_sys_TEA_f0_sop;                                         // Start of packet indicator
logic           usb_sub_sys_TEA_f0_eop;                                         // End of packet indicator
logic    [35:0] usb_sub_sys_TEA_f0_flitdata;                                    // Flit data
logic           usb_sub_sys_TEA_f0_ready;                                       // Flit transfer ready
logic           usb_sub_sys_TEA_f1_activity;                                    // Upcoming activity indicator
logic           usb_sub_sys_TEA_f1_req;                                         // Flit transfer request
logic           usb_sub_sys_TEA_f1_sop;                                         // Start of packet indicator
logic           usb_sub_sys_TEA_f1_eop;                                         // End of packet indicator
logic    [59:0] usb_sub_sys_TEA_f1_flitdata;                                    // Flit data
logic           usb_sub_sys_TEA_f1_ready;                                       // Flit transfer ready
logic           pam3_sub_sys_TEA_f0_activity;                                   // Upcoming activity indicator
logic           pam3_sub_sys_TEA_f0_req;                                        // Flit transfer request
logic           pam3_sub_sys_TEA_f0_sop;                                        // Start of packet indicator
logic           pam3_sub_sys_TEA_f0_eop;                                        // End of packet indicator
logic    [35:0] pam3_sub_sys_TEA_f0_flitdata;                                   // Flit data
logic           pam3_sub_sys_TEA_f0_ready;                                      // Flit transfer ready
logic           pam3_sub_sys_TEA_f1_activity;                                   // Upcoming activity indicator
logic           pam3_sub_sys_TEA_f1_req;                                        // Flit transfer request
logic           pam3_sub_sys_TEA_f1_sop;                                        // Start of packet indicator
logic           pam3_sub_sys_TEA_f1_eop;                                        // End of packet indicator
logic    [59:0] pam3_sub_sys_TEA_f1_flitdata;                                   // Flit data
logic           pam3_sub_sys_TEA_f1_ready;                                      // Flit transfer ready
logic           usb4_phy_TEA_f0_activity;                                       // Upcoming activity indicator
logic           usb4_phy_TEA_f0_req;                                            // Flit transfer request
logic           usb4_phy_TEA_f0_sop;                                            // Start of packet indicator
logic           usb4_phy_TEA_f0_eop;                                            // End of packet indicator
logic    [35:0] usb4_phy_TEA_f0_flitdata;                                       // Flit data
logic           usb4_phy_TEA_f0_ready;                                          // Flit transfer ready
logic           usb4_phy_TEA_f1_activity;                                       // Upcoming activity indicator
logic           usb4_phy_TEA_f1_req;                                            // Flit transfer request
logic           usb4_phy_TEA_f1_sop;                                            // Start of packet indicator
logic           usb4_phy_TEA_f1_eop;                                            // End of packet indicator
logic    [59:0] usb4_phy_TEA_f1_flitdata;                                       // Flit data
logic           usb4_phy_TEA_f1_ready;                                          // Flit transfer ready
logic           pam3_xcvr_TEA_f0_activity;                                      // Upcoming activity indicator
logic           pam3_xcvr_TEA_f0_req;                                           // Flit transfer request
logic           pam3_xcvr_TEA_f0_sop;                                           // Start of packet indicator
logic           pam3_xcvr_TEA_f0_eop;                                           // End of packet indicator
logic    [35:0] pam3_xcvr_TEA_f0_flitdata;                                      // Flit data
logic           pam3_xcvr_TEA_f0_ready;                                         // Flit transfer ready
logic           pam3_xcvr_TEA_f1_activity;                                      // Upcoming activity indicator
logic           pam3_xcvr_TEA_f1_req;                                           // Flit transfer request
logic           pam3_xcvr_TEA_f1_sop;                                           // Start of packet indicator
logic           pam3_xcvr_TEA_f1_eop;                                           // End of packet indicator
logic    [59:0] pam3_xcvr_TEA_f1_flitdata;                                      // Flit data
logic           pam3_xcvr_TEA_f1_ready;                                         // Flit transfer ready
logic           tap2apb_pclk_sync_rst_n;
logic           noc_clk_sync_rst_n;
// param u8            axi4IeaCnt      desc(Count of AXI4-IEA instances);
// param nocAxi4IeaCfg axi4IeaList[1]  desc(List of AXI4-IEA instance configurations);
// param u8            axi4TeaCnt      desc(Count of AXI4-TEA instances);
// param nocAxi4TeaCfg axi4TeaList[1]  desc(List of AXI4-TEA instance configurations);
// param u8            apbIeaCnt       desc(Count of APB-IEA instances);
// param nocApbIeaCfg  apbIeaList[64]  desc(List of APB-IEA instance configurations);
// param u8            apbTeaCnt       desc(Count of APB-TEA instances);
// param nocApbTeaCfg  apbTeaList[64]  desc(List of APB-TEA instance configurations);
// param u8            ahbIeaCnt       desc(Count of AHB-IEA instances);
// param nocAhbIeaCfg  ahbIeaList[64]  desc(List of AHB-IEA instance configurations);
// param u8            ahbTeaCnt       desc(Count of AHB-TEA instances);
// param nocAhbTeaCfg  ahbTeaList[64]  desc(List of AHB-TEA instance configurations);
// param u8                 testNocIOIeaCnt       desc(Count of TESTNOC-IEA instances);
// param testNocIOIeaCfg    testNocIOIeaList[64]  desc(List of TESTNOC-IEA instance configurations);
// param u8                 testNocIOTeaCnt       desc(Count of TESTNOC-TEA instances);
// param testNocIOTeaCfg    testNocIOTeaList[64]  desc(List of TESTNOC-TEA instance configurations);
// param u8            llkpCnt         desc(Count of LLKP instances);
// param nocLlkpCfg    llkpList[64]    desc(List of LLKP instance configurations);
// param u8            lkpCnt          desc(Count of LKP instances);
// param nocLkpCfg     lkpList[64]     desc(List of LKP instance configurations);
// param u8            linkSrcCnt      desc(Count of LINKSRC instances);
// param nocLinkSrcCfg linkSrcList[64] desc(List of LINKSRC instance configurations);
// param u8            linkTgtCnt      desc(Count of LINKTGT instances);
// param nocLinkTgtCfg linkTgtList[64] desc(List of LINKTGT instance configurations);
// param u8            linkCnt         desc(Count of LINK instances);
// param nocLinkCfg    linkList[64]    desc(List of LINK instance configurations);
// param u8            rtrCnt          desc(Count of RTR instances);
// param nocRtrCfg     rtrList[64]     desc(List of RTR instance configurations);
// ============================================
// Clocks and reset
// ============================================
// Loop for each clock source
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// AXI4 Initiator Ports (AXI4 subordinate)
// ============================================
// ============================================
// APB Initiator Ports (APB subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// AHB Initiator Ports (AHB subordinate)
// ============================================
// ============================================
// AXI4 Target Ports (AXI4 manager)
// ============================================
// ============================================
// APB Target Ports (APB manager(s))
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// AHB Target Ports (AHB manager(s))
// ============================================
// ===========================================
// Full Reset Synchronizers (1 for each reset domain)
// ===========================================
usb4_tc_noc_rstFStap2apb_pclk rstFStap2apb_pclk (
  .clk(tap2apb_pclk),                                                           // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(tap2apb_pclk_sync_rst_n),                                          // o:1
  .logicReset()                                                                 // o:1
);
usb4_tc_noc_rstFSnoc_clk rstFSnoc_clk (
  .clk(noc_clk),                                                                // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(noc_clk_sync_rst_n),                                               // o:1
  .logicReset()                                                                 // o:1
);
// ===========================================
// AXI4-IEA Instances
// ===========================================
// ===========================================
// AXI4-TEA Instances
// ===========================================
// ===========================================
// APB-IEA Instances
// ===========================================
usb4_tc_noc_apbiea0 apbiea0 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .s_paddr(apb_mstr_paddr),                                                     // i:32
  .s_psel(apb_mstr_psel),                                                       // i:1
  .s_penable(apb_mstr_penable),                                                 // i:1
  .s_pwrite(apb_mstr_pwrite),                                                   // i:1
  .s_pwdata(apb_mstr_pwdata),                                                   // i:32
  .s_pstrb(apb_mstr_pstrb),                                                     // i:4
  .s_pready(apb_mstr_pready),                                                   // o:1
  .s_prdata(apb_mstr_prdata),                                                   // o:32
  .s_pslverr(apb_mstr_pslverr),                                                 // o:1
  .f0_activity(apb_mstr_f0_activity),                                           // o:1
  .f0_req(apb_mstr_f0_req),                                                     // o:1
  .f0_sop(apb_mstr_f0_sop),                                                     // o:1
  .f0_eop(apb_mstr_f0_eop),                                                     // o:1
  .f0_flitdata(apb_mstr_f0_flitdata),                                           // o:36
  .f0_ready(apb_mstr_f0_ready),                                                 // i:1
  .f1_activity(apb_mstr_f1_activity),                                           // o:1
  .f1_req(apb_mstr_f1_req),                                                     // o:1
  .f1_sop(apb_mstr_f1_sop),                                                     // o:1
  .f1_eop(apb_mstr_f1_eop),                                                     // o:1
  .f1_flitdata(apb_mstr_f1_flitdata),                                           // o:60
  .f1_ready(apb_mstr_f1_ready),                                                 // i:1
  .r0_activity(apb_mstr_r0_activity),                                           // i:1
  .r0_req(apb_mstr_r0_req),                                                     // i:1
  .r0_sop(apb_mstr_r0_sop),                                                     // i:1
  .r0_eop(apb_mstr_r0_eop),                                                     // i:1
  .r0_flitdata(apb_mstr_r0_flitdata),                                           // i:34
  .r0_ready(apb_mstr_r0_ready),                                                 // o:1
  .r1_activity(apb_mstr_r1_activity),                                           // i:1
  .r1_req(apb_mstr_r1_req),                                                     // i:1
  .r1_sop(apb_mstr_r1_sop),                                                     // i:1
  .r1_eop(apb_mstr_r1_eop),                                                     // i:1
  .r1_flitdata(apb_mstr_r1_flitdata),                                           // i:24
  .r1_ready(apb_mstr_r1_ready)                                                  // o:1
);
usb4_tc_noc_apbiea1 apbiea1 (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(tap2apb_pclk_sync_rst_n),                                              // i:1
  .s_paddr(cdb_paddr),                                                          // i:32
  .s_psel(cdb_psel),                                                            // i:1
  .s_penable(cdb_penable),                                                      // i:1
  .s_pwrite(cdb_pwrite),                                                        // i:1
  .s_pwdata(cdb_pwdata),                                                        // i:32
  .s_pstrb(cdb_pstrb),                                                          // i:4
  .s_pready(cdb_pready),                                                        // o:1
  .s_prdata(cdb_prdata),                                                        // o:32
  .s_pslverr(cdb_pslverr),                                                      // o:1
  .f0_activity(tap2apb_f0_activity),                                            // o:1
  .f0_req(tap2apb_f0_req),                                                      // o:1
  .f0_sop(tap2apb_f0_sop),                                                      // o:1
  .f0_eop(tap2apb_f0_eop),                                                      // o:1
  .f0_flitdata(tap2apb_f0_flitdata),                                            // o:36
  .f0_ready(tap2apb_f0_ready),                                                  // i:1
  .f1_activity(tap2apb_f1_activity),                                            // o:1
  .f1_req(tap2apb_f1_req),                                                      // o:1
  .f1_sop(tap2apb_f1_sop),                                                      // o:1
  .f1_eop(tap2apb_f1_eop),                                                      // o:1
  .f1_flitdata(tap2apb_f1_flitdata),                                            // o:60
  .f1_ready(tap2apb_f1_ready),                                                  // i:1
  .r0_activity(tap2apb_r0_activity),                                            // i:1
  .r0_req(tap2apb_r0_req),                                                      // i:1
  .r0_sop(tap2apb_r0_sop),                                                      // i:1
  .r0_eop(tap2apb_r0_eop),                                                      // i:1
  .r0_flitdata(tap2apb_r0_flitdata),                                            // i:34
  .r0_ready(tap2apb_r0_ready),                                                  // o:1
  .r1_activity(tap2apb_r1_activity),                                            // i:1
  .r1_req(tap2apb_r1_req),                                                      // i:1
  .r1_sop(tap2apb_r1_sop),                                                      // i:1
  .r1_eop(tap2apb_r1_eop),                                                      // i:1
  .r1_flitdata(tap2apb_r1_flitdata),                                            // i:24
  .r1_ready(tap2apb_r1_ready)                                                   // o:1
);
// ===========================================
// AHB-IEA Instances
// ===========================================
// ===========================================
// APB-TEA Instances
// ===========================================
usb4_tc_noc_apbtea0 apbtea0 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .t_paddr(cmn_cdb_paddr),                                                      // o:9
  .t_psel(cmn_cdb_psel),                                                        // o:1
  .t_penable(cmn_cdb_penable),                                                  // o:1
  .t_pwrite(cmn_cdb_pwrite),                                                    // o:1
  .t_pwdata(cmn_cdb_pwdata),                                                    // o:32
  .t_pstrb(cmn_cdb_pstrb),                                                      // o:4
  .t_pready(cmn_cdb_pready),                                                    // i:1
  .t_prdata(cmn_cdb_prdata),                                                    // i:32
  .f0_activity(pam3_cmn_TEA_f0_activity),                                       // i:1
  .f0_req(pam3_cmn_TEA_f0_req),                                                 // i:1
  .f0_sop(pam3_cmn_TEA_f0_sop),                                                 // i:1
  .f0_eop(pam3_cmn_TEA_f0_eop),                                                 // i:1
  .f0_flitdata(pam3_cmn_TEA_f0_flitdata),                                       // i:36
  .f0_ready(pam3_cmn_TEA_f0_ready),                                             // o:1
  .f1_activity(pam3_cmn_TEA_f1_activity),                                       // i:1
  .f1_req(pam3_cmn_TEA_f1_req),                                                 // i:1
  .f1_sop(pam3_cmn_TEA_f1_sop),                                                 // i:1
  .f1_eop(pam3_cmn_TEA_f1_eop),                                                 // i:1
  .f1_flitdata(pam3_cmn_TEA_f1_flitdata),                                       // i:60
  .f1_ready(pam3_cmn_TEA_f1_ready),                                             // o:1
  .r0_activity(pam3_cmn_TEA_r0_activity),                                       // o:1
  .r0_req(pam3_cmn_TEA_r0_req),                                                 // o:1
  .r0_sop(pam3_cmn_TEA_r0_sop),                                                 // o:1
  .r0_eop(pam3_cmn_TEA_r0_eop),                                                 // o:1
  .r0_flitdata(pam3_cmn_TEA_r0_flitdata),                                       // o:34
  .r0_ready(pam3_cmn_TEA_r0_ready),                                             // i:1
  .r1_activity(pam3_cmn_TEA_r1_activity),                                       // o:1
  .r1_req(pam3_cmn_TEA_r1_req),                                                 // o:1
  .r1_sop(pam3_cmn_TEA_r1_sop),                                                 // o:1
  .r1_eop(pam3_cmn_TEA_r1_eop),                                                 // o:1
  .r1_flitdata(pam3_cmn_TEA_r1_flitdata),                                       // o:24
  .r1_ready(pam3_cmn_TEA_r1_ready)                                              // i:1
);
usb4_tc_noc_apbtea1 apbtea1 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .t_paddr(tc_reg_paddr),                                                       // o:16
  .t_psel(tc_reg_psel),                                                         // o:1
  .t_penable(tc_reg_penable),                                                   // o:1
  .t_pwrite(tc_reg_pwrite),                                                     // o:1
  .t_pwdata(tc_reg_pwdata),                                                     // o:32
  .t_pstrb(tc_reg_pstrb),                                                       // o:4
  .t_pready(tc_reg_pready),                                                     // i:1
  .t_prdata(tc_reg_prdata),                                                     // i:32
  .f0_activity(tc_reg_TEA_f0_activity),                                         // i:1
  .f0_req(tc_reg_TEA_f0_req),                                                   // i:1
  .f0_sop(tc_reg_TEA_f0_sop),                                                   // i:1
  .f0_eop(tc_reg_TEA_f0_eop),                                                   // i:1
  .f0_flitdata(tc_reg_TEA_f0_flitdata),                                         // i:36
  .f0_ready(tc_reg_TEA_f0_ready),                                               // o:1
  .f1_activity(tc_reg_TEA_f1_activity),                                         // i:1
  .f1_req(tc_reg_TEA_f1_req),                                                   // i:1
  .f1_sop(tc_reg_TEA_f1_sop),                                                   // i:1
  .f1_eop(tc_reg_TEA_f1_eop),                                                   // i:1
  .f1_flitdata(tc_reg_TEA_f1_flitdata),                                         // i:60
  .f1_ready(tc_reg_TEA_f1_ready),                                               // o:1
  .r0_activity(tc_reg_TEA_r0_activity),                                         // o:1
  .r0_req(tc_reg_TEA_r0_req),                                                   // o:1
  .r0_sop(tc_reg_TEA_r0_sop),                                                   // o:1
  .r0_eop(tc_reg_TEA_r0_eop),                                                   // o:1
  .r0_flitdata(tc_reg_TEA_r0_flitdata),                                         // o:34
  .r0_ready(tc_reg_TEA_r0_ready),                                               // i:1
  .r1_activity(tc_reg_TEA_r1_activity),                                         // o:1
  .r1_req(tc_reg_TEA_r1_req),                                                   // o:1
  .r1_sop(tc_reg_TEA_r1_sop),                                                   // o:1
  .r1_eop(tc_reg_TEA_r1_eop),                                                   // o:1
  .r1_flitdata(tc_reg_TEA_r1_flitdata),                                         // o:24
  .r1_ready(tc_reg_TEA_r1_ready)                                                // i:1
);
usb4_tc_noc_apbtea2 apbtea2 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .t_paddr(usb_sub_sys_paddr),                                                  // o:16
  .t_psel(usb_sub_sys_psel),                                                    // o:1
  .t_penable(usb_sub_sys_penable),                                              // o:1
  .t_pwrite(usb_sub_sys_pwrite),                                                // o:1
  .t_pwdata(usb_sub_sys_pwdata),                                                // o:32
  .t_pstrb(usb_sub_sys_pstrb),                                                  // o:4
  .t_pready(usb_sub_sys_pready),                                                // i:1
  .t_prdata(usb_sub_sys_prdata),                                                // i:32
  .f0_activity(usb_sub_sys_TEA_f0_activity),                                    // i:1
  .f0_req(usb_sub_sys_TEA_f0_req),                                              // i:1
  .f0_sop(usb_sub_sys_TEA_f0_sop),                                              // i:1
  .f0_eop(usb_sub_sys_TEA_f0_eop),                                              // i:1
  .f0_flitdata(usb_sub_sys_TEA_f0_flitdata),                                    // i:36
  .f0_ready(usb_sub_sys_TEA_f0_ready),                                          // o:1
  .f1_activity(usb_sub_sys_TEA_f1_activity),                                    // i:1
  .f1_req(usb_sub_sys_TEA_f1_req),                                              // i:1
  .f1_sop(usb_sub_sys_TEA_f1_sop),                                              // i:1
  .f1_eop(usb_sub_sys_TEA_f1_eop),                                              // i:1
  .f1_flitdata(usb_sub_sys_TEA_f1_flitdata),                                    // i:60
  .f1_ready(usb_sub_sys_TEA_f1_ready),                                          // o:1
  .r0_activity(usb_sub_sys_TEA_r0_activity),                                    // o:1
  .r0_req(usb_sub_sys_TEA_r0_req),                                              // o:1
  .r0_sop(usb_sub_sys_TEA_r0_sop),                                              // o:1
  .r0_eop(usb_sub_sys_TEA_r0_eop),                                              // o:1
  .r0_flitdata(usb_sub_sys_TEA_r0_flitdata),                                    // o:34
  .r0_ready(usb_sub_sys_TEA_r0_ready),                                          // i:1
  .r1_activity(usb_sub_sys_TEA_r1_activity),                                    // o:1
  .r1_req(usb_sub_sys_TEA_r1_req),                                              // o:1
  .r1_sop(usb_sub_sys_TEA_r1_sop),                                              // o:1
  .r1_eop(usb_sub_sys_TEA_r1_eop),                                              // o:1
  .r1_flitdata(usb_sub_sys_TEA_r1_flitdata),                                    // o:24
  .r1_ready(usb_sub_sys_TEA_r1_ready)                                           // i:1
);
usb4_tc_noc_apbtea3 apbtea3 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .t_paddr(pam3_sub_sys_paddr),                                                 // o:16
  .t_psel(pam3_sub_sys_psel),                                                   // o:1
  .t_penable(pam3_sub_sys_penable),                                             // o:1
  .t_pwrite(pam3_sub_sys_pwrite),                                               // o:1
  .t_pwdata(pam3_sub_sys_pwdata),                                               // o:32
  .t_pstrb(pam3_sub_sys_pstrb),                                                 // o:4
  .t_pready(pam3_sub_sys_pready),                                               // i:1
  .t_prdata(pam3_sub_sys_prdata),                                               // i:32
  .f0_activity(pam3_sub_sys_TEA_f0_activity),                                   // i:1
  .f0_req(pam3_sub_sys_TEA_f0_req),                                             // i:1
  .f0_sop(pam3_sub_sys_TEA_f0_sop),                                             // i:1
  .f0_eop(pam3_sub_sys_TEA_f0_eop),                                             // i:1
  .f0_flitdata(pam3_sub_sys_TEA_f0_flitdata),                                   // i:36
  .f0_ready(pam3_sub_sys_TEA_f0_ready),                                         // o:1
  .f1_activity(pam3_sub_sys_TEA_f1_activity),                                   // i:1
  .f1_req(pam3_sub_sys_TEA_f1_req),                                             // i:1
  .f1_sop(pam3_sub_sys_TEA_f1_sop),                                             // i:1
  .f1_eop(pam3_sub_sys_TEA_f1_eop),                                             // i:1
  .f1_flitdata(pam3_sub_sys_TEA_f1_flitdata),                                   // i:60
  .f1_ready(pam3_sub_sys_TEA_f1_ready),                                         // o:1
  .r0_activity(pam3_sub_sys_TEA_r0_activity),                                   // o:1
  .r0_req(pam3_sub_sys_TEA_r0_req),                                             // o:1
  .r0_sop(pam3_sub_sys_TEA_r0_sop),                                             // o:1
  .r0_eop(pam3_sub_sys_TEA_r0_eop),                                             // o:1
  .r0_flitdata(pam3_sub_sys_TEA_r0_flitdata),                                   // o:34
  .r0_ready(pam3_sub_sys_TEA_r0_ready),                                         // i:1
  .r1_activity(pam3_sub_sys_TEA_r1_activity),                                   // o:1
  .r1_req(pam3_sub_sys_TEA_r1_req),                                             // o:1
  .r1_sop(pam3_sub_sys_TEA_r1_sop),                                             // o:1
  .r1_eop(pam3_sub_sys_TEA_r1_eop),                                             // o:1
  .r1_flitdata(pam3_sub_sys_TEA_r1_flitdata),                                   // o:24
  .r1_ready(pam3_sub_sys_TEA_r1_ready)                                          // i:1
);
usb4_tc_noc_apbtea4 apbtea4 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .t_paddr(apb_tgt_paddr),                                                      // o:18
  .t_psel(apb_tgt_psel),                                                        // o:1
  .t_penable(apb_tgt_penable),                                                  // o:1
  .t_pwrite(apb_tgt_pwrite),                                                    // o:1
  .t_pwdata(apb_tgt_pwdata),                                                    // o:32
  .t_pstrb(apb_tgt_pstrb),                                                      // o:4
  .t_pready(apb_tgt_pready),                                                    // i:1
  .t_prdata(apb_tgt_prdata),                                                    // i:32
  .t_pslverr(apb_tgt_pslverr),                                                  // i:1
  .f0_activity(usb4_phy_TEA_f0_activity),                                       // i:1
  .f0_req(usb4_phy_TEA_f0_req),                                                 // i:1
  .f0_sop(usb4_phy_TEA_f0_sop),                                                 // i:1
  .f0_eop(usb4_phy_TEA_f0_eop),                                                 // i:1
  .f0_flitdata(usb4_phy_TEA_f0_flitdata),                                       // i:36
  .f0_ready(usb4_phy_TEA_f0_ready),                                             // o:1
  .f1_activity(usb4_phy_TEA_f1_activity),                                       // i:1
  .f1_req(usb4_phy_TEA_f1_req),                                                 // i:1
  .f1_sop(usb4_phy_TEA_f1_sop),                                                 // i:1
  .f1_eop(usb4_phy_TEA_f1_eop),                                                 // i:1
  .f1_flitdata(usb4_phy_TEA_f1_flitdata),                                       // i:60
  .f1_ready(usb4_phy_TEA_f1_ready),                                             // o:1
  .r0_activity(usb4_phy_TEA_r0_activity),                                       // o:1
  .r0_req(usb4_phy_TEA_r0_req),                                                 // o:1
  .r0_sop(usb4_phy_TEA_r0_sop),                                                 // o:1
  .r0_eop(usb4_phy_TEA_r0_eop),                                                 // o:1
  .r0_flitdata(usb4_phy_TEA_r0_flitdata),                                       // o:34
  .r0_ready(usb4_phy_TEA_r0_ready),                                             // i:1
  .r1_activity(usb4_phy_TEA_r1_activity),                                       // o:1
  .r1_req(usb4_phy_TEA_r1_req),                                                 // o:1
  .r1_sop(usb4_phy_TEA_r1_sop),                                                 // o:1
  .r1_eop(usb4_phy_TEA_r1_eop),                                                 // o:1
  .r1_flitdata(usb4_phy_TEA_r1_flitdata),                                       // o:24
  .r1_ready(usb4_phy_TEA_r1_ready)                                              // i:1
);
usb4_tc_noc_apbtea5 apbtea5 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .t_paddr(xcvr_ln_0_paddr),                                                    // o:10
  .t_psel(xcvr_ln_0_psel),                                                      // o:1
  .t_penable(xcvr_ln_0_penable),                                                // o:1
  .t_pwrite(xcvr_ln_0_pwrite),                                                  // o:1
  .t_pwdata(xcvr_ln_0_pwdata),                                                  // o:32
  .t_pstrb(xcvr_ln_0_pstrb),                                                    // o:4
  .t_pready(xcvr_ln_0_pready),                                                  // i:1
  .t_prdata(xcvr_ln_0_prdata),                                                  // i:32
  .f0_activity(pam3_xcvr_TEA_f0_activity),                                      // i:1
  .f0_req(pam3_xcvr_TEA_f0_req),                                                // i:1
  .f0_sop(pam3_xcvr_TEA_f0_sop),                                                // i:1
  .f0_eop(pam3_xcvr_TEA_f0_eop),                                                // i:1
  .f0_flitdata(pam3_xcvr_TEA_f0_flitdata),                                      // i:36
  .f0_ready(pam3_xcvr_TEA_f0_ready),                                            // o:1
  .f1_activity(pam3_xcvr_TEA_f1_activity),                                      // i:1
  .f1_req(pam3_xcvr_TEA_f1_req),                                                // i:1
  .f1_sop(pam3_xcvr_TEA_f1_sop),                                                // i:1
  .f1_eop(pam3_xcvr_TEA_f1_eop),                                                // i:1
  .f1_flitdata(pam3_xcvr_TEA_f1_flitdata),                                      // i:60
  .f1_ready(pam3_xcvr_TEA_f1_ready),                                            // o:1
  .r0_activity(pam3_xcvr_TEA_r0_activity),                                      // o:1
  .r0_req(pam3_xcvr_TEA_r0_req),                                                // o:1
  .r0_sop(pam3_xcvr_TEA_r0_sop),                                                // o:1
  .r0_eop(pam3_xcvr_TEA_r0_eop),                                                // o:1
  .r0_flitdata(pam3_xcvr_TEA_r0_flitdata),                                      // o:34
  .r0_ready(pam3_xcvr_TEA_r0_ready),                                            // i:1
  .r1_activity(pam3_xcvr_TEA_r1_activity),                                      // o:1
  .r1_req(pam3_xcvr_TEA_r1_req),                                                // o:1
  .r1_sop(pam3_xcvr_TEA_r1_sop),                                                // o:1
  .r1_eop(pam3_xcvr_TEA_r1_eop),                                                // o:1
  .r1_flitdata(pam3_xcvr_TEA_r1_flitdata),                                      // o:24
  .r1_ready(pam3_xcvr_TEA_r1_ready)                                             // i:1
);
// ===========================================
// AHB-TEA Instances
// ===========================================
// ===========================================
// Link Instances
// ===========================================
usb4_tc_noc_link0 link0 (
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .slf0_activity(tap2apb_f0_activity),                                          // i:1
  .slf0_req(tap2apb_f0_req),                                                    // i:1
  .slf0_sop(tap2apb_f0_sop),                                                    // i:1
  .slf0_eop(tap2apb_f0_eop),                                                    // i:1
  .slf0_flitdata(tap2apb_f0_flitdata),                                          // i:36
  .slf0_ready(tap2apb_f0_ready),                                                // o:1
  .slf1_activity(tap2apb_f1_activity),                                          // i:1
  .slf1_req(tap2apb_f1_req),                                                    // i:1
  .slf1_sop(tap2apb_f1_sop),                                                    // i:1
  .slf1_eop(tap2apb_f1_eop),                                                    // i:1
  .slf1_flitdata(tap2apb_f1_flitdata),                                          // i:60
  .slf1_ready(tap2apb_f1_ready),                                                // o:1
  .slr0_activity(tap2apb_r0_activity),                                          // o:1
  .slr0_req(tap2apb_r0_req),                                                    // o:1
  .slr0_sop(tap2apb_r0_sop),                                                    // o:1
  .slr0_eop(tap2apb_r0_eop),                                                    // o:1
  .slr0_flitdata(tap2apb_r0_flitdata),                                          // o:34
  .slr0_ready(tap2apb_r0_ready),                                                // i:1
  .slr1_activity(tap2apb_r1_activity),                                          // o:1
  .slr1_req(tap2apb_r1_req),                                                    // o:1
  .slr1_sop(tap2apb_r1_sop),                                                    // o:1
  .slr1_eop(tap2apb_r1_eop),                                                    // o:1
  .slr1_flitdata(tap2apb_r1_flitdata),                                          // o:24
  .slr1_ready(tap2apb_r1_ready),                                                // i:1
  .dlf0_activity(RTR_INI0_f0_activity),                                         // o:1
  .dlf0_req(RTR_INI0_f0_req),                                                   // o:1
  .dlf0_sop(RTR_INI0_f0_sop),                                                   // o:1
  .dlf0_eop(RTR_INI0_f0_eop),                                                   // o:1
  .dlf0_flitdata(RTR_INI0_f0_flitdata),                                         // o:36
  .dlf0_ready(RTR_INI0_f0_ready),                                               // i:1
  .dlf1_activity(RTR_INI0_f1_activity),                                         // o:1
  .dlf1_req(RTR_INI0_f1_req),                                                   // o:1
  .dlf1_sop(RTR_INI0_f1_sop),                                                   // o:1
  .dlf1_eop(RTR_INI0_f1_eop),                                                   // o:1
  .dlf1_flitdata(RTR_INI0_f1_flitdata),                                         // o:60
  .dlf1_ready(RTR_INI0_f1_ready),                                               // i:1
  .dlr0_activity(RTR_INI0_r0_activity),                                         // i:1
  .dlr0_req(RTR_INI0_r0_req),                                                   // i:1
  .dlr0_sop(RTR_INI0_r0_sop),                                                   // i:1
  .dlr0_eop(RTR_INI0_r0_eop),                                                   // i:1
  .dlr0_flitdata(RTR_INI0_r0_flitdata),                                         // i:34
  .dlr0_ready(RTR_INI0_r0_ready),                                               // o:1
  .dlr1_activity(RTR_INI0_r1_activity),                                         // i:1
  .dlr1_req(RTR_INI0_r1_req),                                                   // i:1
  .dlr1_sop(RTR_INI0_r1_sop),                                                   // i:1
  .dlr1_eop(RTR_INI0_r1_eop),                                                   // i:1
  .dlr1_flitdata(RTR_INI0_r1_flitdata),                                         // i:24
  .dlr1_ready(RTR_INI0_r1_ready)                                                // o:1
);
// ===========================================
// LLink Instances
// ===========================================
// ===========================================
// Router Instances
// ===========================================
usb4_tc_noc_rtr0 rtr0 (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .apb_mstr_f0_activity(apb_mstr_f0_activity),                                  // i:1
  .apb_mstr_f0_req(apb_mstr_f0_req),                                            // i:1
  .apb_mstr_f0_sop(apb_mstr_f0_sop),                                            // i:1
  .apb_mstr_f0_eop(apb_mstr_f0_eop),                                            // i:1
  .apb_mstr_f0_flitdata(apb_mstr_f0_flitdata),                                  // i:36
  .apb_mstr_f0_ready(apb_mstr_f0_ready),                                        // o:1
  .apb_mstr_f1_activity(apb_mstr_f1_activity),                                  // i:1
  .apb_mstr_f1_req(apb_mstr_f1_req),                                            // i:1
  .apb_mstr_f1_sop(apb_mstr_f1_sop),                                            // i:1
  .apb_mstr_f1_eop(apb_mstr_f1_eop),                                            // i:1
  .apb_mstr_f1_flitdata(apb_mstr_f1_flitdata),                                  // i:60
  .apb_mstr_f1_ready(apb_mstr_f1_ready),                                        // o:1
  .apb_mstr_r0_activity(apb_mstr_r0_activity),                                  // o:1
  .apb_mstr_r0_req(apb_mstr_r0_req),                                            // o:1
  .apb_mstr_r0_sop(apb_mstr_r0_sop),                                            // o:1
  .apb_mstr_r0_eop(apb_mstr_r0_eop),                                            // o:1
  .apb_mstr_r0_flitdata(apb_mstr_r0_flitdata),                                  // o:34
  .apb_mstr_r0_ready(apb_mstr_r0_ready),                                        // i:1
  .apb_mstr_r1_activity(apb_mstr_r1_activity),                                  // o:1
  .apb_mstr_r1_req(apb_mstr_r1_req),                                            // o:1
  .apb_mstr_r1_sop(apb_mstr_r1_sop),                                            // o:1
  .apb_mstr_r1_eop(apb_mstr_r1_eop),                                            // o:1
  .apb_mstr_r1_flitdata(apb_mstr_r1_flitdata),                                  // o:24
  .apb_mstr_r1_ready(apb_mstr_r1_ready),                                        // i:1
  .RTR_INI0_f0_activity(RTR_INI0_f0_activity),                                  // i:1
  .RTR_INI0_f0_req(RTR_INI0_f0_req),                                            // i:1
  .RTR_INI0_f0_sop(RTR_INI0_f0_sop),                                            // i:1
  .RTR_INI0_f0_eop(RTR_INI0_f0_eop),                                            // i:1
  .RTR_INI0_f0_flitdata(RTR_INI0_f0_flitdata),                                  // i:36
  .RTR_INI0_f0_ready(RTR_INI0_f0_ready),                                        // o:1
  .RTR_INI0_f1_activity(RTR_INI0_f1_activity),                                  // i:1
  .RTR_INI0_f1_req(RTR_INI0_f1_req),                                            // i:1
  .RTR_INI0_f1_sop(RTR_INI0_f1_sop),                                            // i:1
  .RTR_INI0_f1_eop(RTR_INI0_f1_eop),                                            // i:1
  .RTR_INI0_f1_flitdata(RTR_INI0_f1_flitdata),                                  // i:60
  .RTR_INI0_f1_ready(RTR_INI0_f1_ready),                                        // o:1
  .RTR_INI0_r0_activity(RTR_INI0_r0_activity),                                  // o:1
  .RTR_INI0_r0_req(RTR_INI0_r0_req),                                            // o:1
  .RTR_INI0_r0_sop(RTR_INI0_r0_sop),                                            // o:1
  .RTR_INI0_r0_eop(RTR_INI0_r0_eop),                                            // o:1
  .RTR_INI0_r0_flitdata(RTR_INI0_r0_flitdata),                                  // o:34
  .RTR_INI0_r0_ready(RTR_INI0_r0_ready),                                        // i:1
  .RTR_INI0_r1_activity(RTR_INI0_r1_activity),                                  // o:1
  .RTR_INI0_r1_req(RTR_INI0_r1_req),                                            // o:1
  .RTR_INI0_r1_sop(RTR_INI0_r1_sop),                                            // o:1
  .RTR_INI0_r1_eop(RTR_INI0_r1_eop),                                            // o:1
  .RTR_INI0_r1_flitdata(RTR_INI0_r1_flitdata),                                  // o:24
  .RTR_INI0_r1_ready(RTR_INI0_r1_ready),                                        // i:1
  .pam3_cmn_TEA_f0_activity(pam3_cmn_TEA_f0_activity),                          // o:1
  .pam3_cmn_TEA_f0_req(pam3_cmn_TEA_f0_req),                                    // o:1
  .pam3_cmn_TEA_f0_sop(pam3_cmn_TEA_f0_sop),                                    // o:1
  .pam3_cmn_TEA_f0_eop(pam3_cmn_TEA_f0_eop),                                    // o:1
  .pam3_cmn_TEA_f0_flitdata(pam3_cmn_TEA_f0_flitdata),                          // o:36
  .pam3_cmn_TEA_f0_ready(pam3_cmn_TEA_f0_ready),                                // i:1
  .pam3_cmn_TEA_f1_activity(pam3_cmn_TEA_f1_activity),                          // o:1
  .pam3_cmn_TEA_f1_req(pam3_cmn_TEA_f1_req),                                    // o:1
  .pam3_cmn_TEA_f1_sop(pam3_cmn_TEA_f1_sop),                                    // o:1
  .pam3_cmn_TEA_f1_eop(pam3_cmn_TEA_f1_eop),                                    // o:1
  .pam3_cmn_TEA_f1_flitdata(pam3_cmn_TEA_f1_flitdata),                          // o:60
  .pam3_cmn_TEA_f1_ready(pam3_cmn_TEA_f1_ready),                                // i:1
  .pam3_cmn_TEA_r0_activity(pam3_cmn_TEA_r0_activity),                          // i:1
  .pam3_cmn_TEA_r0_req(pam3_cmn_TEA_r0_req),                                    // i:1
  .pam3_cmn_TEA_r0_sop(pam3_cmn_TEA_r0_sop),                                    // i:1
  .pam3_cmn_TEA_r0_eop(pam3_cmn_TEA_r0_eop),                                    // i:1
  .pam3_cmn_TEA_r0_flitdata(pam3_cmn_TEA_r0_flitdata),                          // i:34
  .pam3_cmn_TEA_r0_ready(pam3_cmn_TEA_r0_ready),                                // o:1
  .pam3_cmn_TEA_r1_activity(pam3_cmn_TEA_r1_activity),                          // i:1
  .pam3_cmn_TEA_r1_req(pam3_cmn_TEA_r1_req),                                    // i:1
  .pam3_cmn_TEA_r1_sop(pam3_cmn_TEA_r1_sop),                                    // i:1
  .pam3_cmn_TEA_r1_eop(pam3_cmn_TEA_r1_eop),                                    // i:1
  .pam3_cmn_TEA_r1_flitdata(pam3_cmn_TEA_r1_flitdata),                          // i:24
  .pam3_cmn_TEA_r1_ready(pam3_cmn_TEA_r1_ready),                                // o:1
  .tc_reg_TEA_f0_activity(tc_reg_TEA_f0_activity),                              // o:1
  .tc_reg_TEA_f0_req(tc_reg_TEA_f0_req),                                        // o:1
  .tc_reg_TEA_f0_sop(tc_reg_TEA_f0_sop),                                        // o:1
  .tc_reg_TEA_f0_eop(tc_reg_TEA_f0_eop),                                        // o:1
  .tc_reg_TEA_f0_flitdata(tc_reg_TEA_f0_flitdata),                              // o:36
  .tc_reg_TEA_f0_ready(tc_reg_TEA_f0_ready),                                    // i:1
  .tc_reg_TEA_f1_activity(tc_reg_TEA_f1_activity),                              // o:1
  .tc_reg_TEA_f1_req(tc_reg_TEA_f1_req),                                        // o:1
  .tc_reg_TEA_f1_sop(tc_reg_TEA_f1_sop),                                        // o:1
  .tc_reg_TEA_f1_eop(tc_reg_TEA_f1_eop),                                        // o:1
  .tc_reg_TEA_f1_flitdata(tc_reg_TEA_f1_flitdata),                              // o:60
  .tc_reg_TEA_f1_ready(tc_reg_TEA_f1_ready),                                    // i:1
  .tc_reg_TEA_r0_activity(tc_reg_TEA_r0_activity),                              // i:1
  .tc_reg_TEA_r0_req(tc_reg_TEA_r0_req),                                        // i:1
  .tc_reg_TEA_r0_sop(tc_reg_TEA_r0_sop),                                        // i:1
  .tc_reg_TEA_r0_eop(tc_reg_TEA_r0_eop),                                        // i:1
  .tc_reg_TEA_r0_flitdata(tc_reg_TEA_r0_flitdata),                              // i:34
  .tc_reg_TEA_r0_ready(tc_reg_TEA_r0_ready),                                    // o:1
  .tc_reg_TEA_r1_activity(tc_reg_TEA_r1_activity),                              // i:1
  .tc_reg_TEA_r1_req(tc_reg_TEA_r1_req),                                        // i:1
  .tc_reg_TEA_r1_sop(tc_reg_TEA_r1_sop),                                        // i:1
  .tc_reg_TEA_r1_eop(tc_reg_TEA_r1_eop),                                        // i:1
  .tc_reg_TEA_r1_flitdata(tc_reg_TEA_r1_flitdata),                              // i:24
  .tc_reg_TEA_r1_ready(tc_reg_TEA_r1_ready),                                    // o:1
  .usb_sub_sys_TEA_f0_activity(usb_sub_sys_TEA_f0_activity),                    // o:1
  .usb_sub_sys_TEA_f0_req(usb_sub_sys_TEA_f0_req),                              // o:1
  .usb_sub_sys_TEA_f0_sop(usb_sub_sys_TEA_f0_sop),                              // o:1
  .usb_sub_sys_TEA_f0_eop(usb_sub_sys_TEA_f0_eop),                              // o:1
  .usb_sub_sys_TEA_f0_flitdata(usb_sub_sys_TEA_f0_flitdata),                    // o:36
  .usb_sub_sys_TEA_f0_ready(usb_sub_sys_TEA_f0_ready),                          // i:1
  .usb_sub_sys_TEA_f1_activity(usb_sub_sys_TEA_f1_activity),                    // o:1
  .usb_sub_sys_TEA_f1_req(usb_sub_sys_TEA_f1_req),                              // o:1
  .usb_sub_sys_TEA_f1_sop(usb_sub_sys_TEA_f1_sop),                              // o:1
  .usb_sub_sys_TEA_f1_eop(usb_sub_sys_TEA_f1_eop),                              // o:1
  .usb_sub_sys_TEA_f1_flitdata(usb_sub_sys_TEA_f1_flitdata),                    // o:60
  .usb_sub_sys_TEA_f1_ready(usb_sub_sys_TEA_f1_ready),                          // i:1
  .usb_sub_sys_TEA_r0_activity(usb_sub_sys_TEA_r0_activity),                    // i:1
  .usb_sub_sys_TEA_r0_req(usb_sub_sys_TEA_r0_req),                              // i:1
  .usb_sub_sys_TEA_r0_sop(usb_sub_sys_TEA_r0_sop),                              // i:1
  .usb_sub_sys_TEA_r0_eop(usb_sub_sys_TEA_r0_eop),                              // i:1
  .usb_sub_sys_TEA_r0_flitdata(usb_sub_sys_TEA_r0_flitdata),                    // i:34
  .usb_sub_sys_TEA_r0_ready(usb_sub_sys_TEA_r0_ready),                          // o:1
  .usb_sub_sys_TEA_r1_activity(usb_sub_sys_TEA_r1_activity),                    // i:1
  .usb_sub_sys_TEA_r1_req(usb_sub_sys_TEA_r1_req),                              // i:1
  .usb_sub_sys_TEA_r1_sop(usb_sub_sys_TEA_r1_sop),                              // i:1
  .usb_sub_sys_TEA_r1_eop(usb_sub_sys_TEA_r1_eop),                              // i:1
  .usb_sub_sys_TEA_r1_flitdata(usb_sub_sys_TEA_r1_flitdata),                    // i:24
  .usb_sub_sys_TEA_r1_ready(usb_sub_sys_TEA_r1_ready),                          // o:1
  .pam3_sub_sys_TEA_f0_activity(pam3_sub_sys_TEA_f0_activity),                  // o:1
  .pam3_sub_sys_TEA_f0_req(pam3_sub_sys_TEA_f0_req),                            // o:1
  .pam3_sub_sys_TEA_f0_sop(pam3_sub_sys_TEA_f0_sop),                            // o:1
  .pam3_sub_sys_TEA_f0_eop(pam3_sub_sys_TEA_f0_eop),                            // o:1
  .pam3_sub_sys_TEA_f0_flitdata(pam3_sub_sys_TEA_f0_flitdata),                  // o:36
  .pam3_sub_sys_TEA_f0_ready(pam3_sub_sys_TEA_f0_ready),                        // i:1
  .pam3_sub_sys_TEA_f1_activity(pam3_sub_sys_TEA_f1_activity),                  // o:1
  .pam3_sub_sys_TEA_f1_req(pam3_sub_sys_TEA_f1_req),                            // o:1
  .pam3_sub_sys_TEA_f1_sop(pam3_sub_sys_TEA_f1_sop),                            // o:1
  .pam3_sub_sys_TEA_f1_eop(pam3_sub_sys_TEA_f1_eop),                            // o:1
  .pam3_sub_sys_TEA_f1_flitdata(pam3_sub_sys_TEA_f1_flitdata),                  // o:60
  .pam3_sub_sys_TEA_f1_ready(pam3_sub_sys_TEA_f1_ready),                        // i:1
  .pam3_sub_sys_TEA_r0_activity(pam3_sub_sys_TEA_r0_activity),                  // i:1
  .pam3_sub_sys_TEA_r0_req(pam3_sub_sys_TEA_r0_req),                            // i:1
  .pam3_sub_sys_TEA_r0_sop(pam3_sub_sys_TEA_r0_sop),                            // i:1
  .pam3_sub_sys_TEA_r0_eop(pam3_sub_sys_TEA_r0_eop),                            // i:1
  .pam3_sub_sys_TEA_r0_flitdata(pam3_sub_sys_TEA_r0_flitdata),                  // i:34
  .pam3_sub_sys_TEA_r0_ready(pam3_sub_sys_TEA_r0_ready),                        // o:1
  .pam3_sub_sys_TEA_r1_activity(pam3_sub_sys_TEA_r1_activity),                  // i:1
  .pam3_sub_sys_TEA_r1_req(pam3_sub_sys_TEA_r1_req),                            // i:1
  .pam3_sub_sys_TEA_r1_sop(pam3_sub_sys_TEA_r1_sop),                            // i:1
  .pam3_sub_sys_TEA_r1_eop(pam3_sub_sys_TEA_r1_eop),                            // i:1
  .pam3_sub_sys_TEA_r1_flitdata(pam3_sub_sys_TEA_r1_flitdata),                  // i:24
  .pam3_sub_sys_TEA_r1_ready(pam3_sub_sys_TEA_r1_ready),                        // o:1
  .usb4_phy_TEA_f0_activity(usb4_phy_TEA_f0_activity),                          // o:1
  .usb4_phy_TEA_f0_req(usb4_phy_TEA_f0_req),                                    // o:1
  .usb4_phy_TEA_f0_sop(usb4_phy_TEA_f0_sop),                                    // o:1
  .usb4_phy_TEA_f0_eop(usb4_phy_TEA_f0_eop),                                    // o:1
  .usb4_phy_TEA_f0_flitdata(usb4_phy_TEA_f0_flitdata),                          // o:36
  .usb4_phy_TEA_f0_ready(usb4_phy_TEA_f0_ready),                                // i:1
  .usb4_phy_TEA_f1_activity(usb4_phy_TEA_f1_activity),                          // o:1
  .usb4_phy_TEA_f1_req(usb4_phy_TEA_f1_req),                                    // o:1
  .usb4_phy_TEA_f1_sop(usb4_phy_TEA_f1_sop),                                    // o:1
  .usb4_phy_TEA_f1_eop(usb4_phy_TEA_f1_eop),                                    // o:1
  .usb4_phy_TEA_f1_flitdata(usb4_phy_TEA_f1_flitdata),                          // o:60
  .usb4_phy_TEA_f1_ready(usb4_phy_TEA_f1_ready),                                // i:1
  .usb4_phy_TEA_r0_activity(usb4_phy_TEA_r0_activity),                          // i:1
  .usb4_phy_TEA_r0_req(usb4_phy_TEA_r0_req),                                    // i:1
  .usb4_phy_TEA_r0_sop(usb4_phy_TEA_r0_sop),                                    // i:1
  .usb4_phy_TEA_r0_eop(usb4_phy_TEA_r0_eop),                                    // i:1
  .usb4_phy_TEA_r0_flitdata(usb4_phy_TEA_r0_flitdata),                          // i:34
  .usb4_phy_TEA_r0_ready(usb4_phy_TEA_r0_ready),                                // o:1
  .usb4_phy_TEA_r1_activity(usb4_phy_TEA_r1_activity),                          // i:1
  .usb4_phy_TEA_r1_req(usb4_phy_TEA_r1_req),                                    // i:1
  .usb4_phy_TEA_r1_sop(usb4_phy_TEA_r1_sop),                                    // i:1
  .usb4_phy_TEA_r1_eop(usb4_phy_TEA_r1_eop),                                    // i:1
  .usb4_phy_TEA_r1_flitdata(usb4_phy_TEA_r1_flitdata),                          // i:24
  .usb4_phy_TEA_r1_ready(usb4_phy_TEA_r1_ready),                                // o:1
  .pam3_xcvr_TEA_f0_activity(pam3_xcvr_TEA_f0_activity),                        // o:1
  .pam3_xcvr_TEA_f0_req(pam3_xcvr_TEA_f0_req),                                  // o:1
  .pam3_xcvr_TEA_f0_sop(pam3_xcvr_TEA_f0_sop),                                  // o:1
  .pam3_xcvr_TEA_f0_eop(pam3_xcvr_TEA_f0_eop),                                  // o:1
  .pam3_xcvr_TEA_f0_flitdata(pam3_xcvr_TEA_f0_flitdata),                        // o:36
  .pam3_xcvr_TEA_f0_ready(pam3_xcvr_TEA_f0_ready),                              // i:1
  .pam3_xcvr_TEA_f1_activity(pam3_xcvr_TEA_f1_activity),                        // o:1
  .pam3_xcvr_TEA_f1_req(pam3_xcvr_TEA_f1_req),                                  // o:1
  .pam3_xcvr_TEA_f1_sop(pam3_xcvr_TEA_f1_sop),                                  // o:1
  .pam3_xcvr_TEA_f1_eop(pam3_xcvr_TEA_f1_eop),                                  // o:1
  .pam3_xcvr_TEA_f1_flitdata(pam3_xcvr_TEA_f1_flitdata),                        // o:60
  .pam3_xcvr_TEA_f1_ready(pam3_xcvr_TEA_f1_ready),                              // i:1
  .pam3_xcvr_TEA_r0_activity(pam3_xcvr_TEA_r0_activity),                        // i:1
  .pam3_xcvr_TEA_r0_req(pam3_xcvr_TEA_r0_req),                                  // i:1
  .pam3_xcvr_TEA_r0_sop(pam3_xcvr_TEA_r0_sop),                                  // i:1
  .pam3_xcvr_TEA_r0_eop(pam3_xcvr_TEA_r0_eop),                                  // i:1
  .pam3_xcvr_TEA_r0_flitdata(pam3_xcvr_TEA_r0_flitdata),                        // i:34
  .pam3_xcvr_TEA_r0_ready(pam3_xcvr_TEA_r0_ready),                              // o:1
  .pam3_xcvr_TEA_r1_activity(pam3_xcvr_TEA_r1_activity),                        // i:1
  .pam3_xcvr_TEA_r1_req(pam3_xcvr_TEA_r1_req),                                  // i:1
  .pam3_xcvr_TEA_r1_sop(pam3_xcvr_TEA_r1_sop),                                  // i:1
  .pam3_xcvr_TEA_r1_eop(pam3_xcvr_TEA_r1_eop),                                  // i:1
  .pam3_xcvr_TEA_r1_flitdata(pam3_xcvr_TEA_r1_flitdata),                        // i:24
  .pam3_xcvr_TEA_r1_ready(pam3_xcvr_TEA_r1_ready)                               // o:1
);
// These coded instructions, statements, and computer programs are the
// copyrighted works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without
// the prior written consent of Cadence Design Systems Inc.
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rstFStap2apb_pclk (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer3 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rstFSnoc_clk (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer3 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0 (
  input  wire            clk,
  input  wire            rst_n,
  // s
  input  wire     [31:0] s_paddr,                                               // Address
  input  wire            s_psel,                                                // Select
  input  wire            s_penable,                                             // Enable
  input  wire            s_pwrite,                                              // Write not read
  input  wire     [31:0] s_pwdata,                                              // Write data
  input  wire      [3:0] s_pstrb,                                               // Write strobes
  output logic           s_pready,                                              // Ready
  output logic    [31:0] s_prdata,                                              // Read data
  output logic           s_pslverr,                                             // Slave error
  // f0
  output logic           f0_activity,                                           // Upcoming activity indicator
  output logic           f0_req,                                                // Flit transfer request
  output logic           f0_sop,                                                // Start of packet indicator
  output logic           f0_eop,                                                // End of packet indicator
  output logic    [35:0] f0_flitdata,                                           // Flit data
  input  wire            f0_ready,                                              // Flit transfer ready
  // f1
  output logic           f1_activity,                                           // Upcoming activity indicator
  output logic           f1_req,                                                // Flit transfer request
  output logic           f1_sop,                                                // Start of packet indicator
  output logic           f1_eop,                                                // End of packet indicator
  output logic    [59:0] f1_flitdata,                                           // Flit data
  input  wire            f1_ready,                                              // Flit transfer ready
  // r0
  input  wire            r0_activity,                                           // Upcoming activity indicator
  input  wire            r0_req,                                                // Flit transfer request
  input  wire            r0_sop,                                                // Start of packet indicator
  input  wire            r0_eop,                                                // End of packet indicator
  input  wire     [33:0] r0_flitdata,                                           // Flit data
  output logic           r0_ready,                                              // Flit transfer ready
  // r1
  input  wire            r1_activity,                                           // Upcoming activity indicator
  input  wire            r1_req,                                                // Flit transfer request
  input  wire            r1_sop,                                                // Start of packet indicator
  input  wire            r1_eop,                                                // End of packet indicator
  input  wire     [23:0] r1_flitdata,                                           // Flit data
  output logic           r1_ready                                               // Flit transfer ready
);

logic    [31:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           int_pslverr;                                                    // Slave error
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic     [2:0] rc_did;
logic     [2:0] rc_sid;
logic    [59:0] rc_hdr;
logic    [31:0] rc_rawAddr;
logic    [31:0] rc_mapdAddr;
logic           rs_buf_we;
logic    [67:0] rs_bus;
logic    [33:0] rds_bus;
logic    [31:0] rds_data;
logic     [1:0] rds_status;
logic     [2:0] wcd_did;
logic     [2:0] wcd_sid;
logic    [71:0] wcd_hdr;
logic    [35:0] wcd_pld;
logic    [31:0] wcd_rawAddr;
logic    [31:0] wcd_mapdAddr;
logic           ws_buf_we;
logic    [23:0] ws_bus;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           gclk;
logic           gclkAct;
logic           gclkEn;
logic     [2:0] rtmp_did;
logic           rtmp_valid;
logic     [2:0] wtmp_did;
logic           wtmp_valid;
logic     [2:0] rpaylen;
logic     [2:0] wpaylen;
logic    [23:0] ws_buf [0:0];
logic     [0:0] ws_buf_en;
logic     [0:0] fcnt;
logic     [0:0] fcnt_nxt;
logic     [0:0] fcnt_en;
logic    [33:0] rs_buf [1:0];
logic     [1:0] rs_buf_en;
logic    [33:0] readSeg;
logic     [2:0] state;
logic     [2:0] state_nxt;
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Initiator Ports (APB subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Ingress APB Pipeline Component
usb4_tc_noc_apbiea0_ipipe ipipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(s_paddr),                                                          // i:32
  .src_psel(s_psel),                                                            // i:1
  .src_penable(s_penable),                                                      // i:1
  .src_pwrite(s_pwrite),                                                        // i:1
  .src_pwdata(s_pwdata),                                                        // i:32
  .src_pstrb(s_pstrb),                                                          // i:4
  .src_pready(s_pready),                                                        // o:1
  .src_prdata(s_prdata),                                                        // o:32
  .src_pslverr(s_pslverr),                                                      // o:1
  .dst_paddr(int_paddr),                                                        // o:32
  .dst_psel(int_psel),                                                          // o:1
  .dst_penable(int_penable),                                                    // o:1
  .dst_pwrite(int_pwrite),                                                      // o:1
  .dst_pwdata(int_pwdata),                                                      // o:32
  .dst_pstrb(int_pstrb),                                                        // o:4
  .dst_pready(int_pready),                                                      // i:1
  .dst_prdata(int_prdata),                                                      // i:32
  .dst_pslverr(int_pslverr)                                                     // i:1
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbiea0_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(if0_activity),                                                  // i:1
  .src_req(if0_req),                                                            // i:1
  .src_sop(if0_sop),                                                            // i:1
  .src_eop(if0_eop),                                                            // i:1
  .src_flitdata(if0_flitdata),                                                  // i:36
  .src_ready(if0_ready),                                                        // o:1
  .dst_activity(f0_activity),                                                   // o:1
  .dst_req(f0_req),                                                             // o:1
  .dst_sop(f0_sop),                                                             // o:1
  .dst_eop(f0_eop),                                                             // o:1
  .dst_flitdata(f0_flitdata),                                                   // o:36
  .dst_ready(f0_ready)                                                          // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbiea0_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(if1_activity),                                                  // i:1
  .src_req(if1_req),                                                            // i:1
  .src_sop(if1_sop),                                                            // i:1
  .src_eop(if1_eop),                                                            // i:1
  .src_flitdata(if1_flitdata),                                                  // i:60
  .src_ready(if1_ready),                                                        // o:1
  .dst_activity(f1_activity),                                                   // o:1
  .dst_req(f1_req),                                                             // o:1
  .dst_sop(f1_sop),                                                             // o:1
  .dst_eop(f1_eop),                                                             // o:1
  .dst_flitdata(f1_flitdata),                                                   // o:60
  .dst_ready(f1_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbiea0_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(r0_activity),                                                   // i:1
  .src_req(r0_req),                                                             // i:1
  .src_sop(r0_sop),                                                             // i:1
  .src_eop(r0_eop),                                                             // i:1
  .src_flitdata(r0_flitdata),                                                   // i:34
  .src_ready(r0_ready),                                                         // o:1
  .dst_activity(ir0_activity),                                                  // o:1
  .dst_req(ir0_req),                                                            // o:1
  .dst_sop(ir0_sop),                                                            // o:1
  .dst_eop(ir0_eop),                                                            // o:1
  .dst_flitdata(ir0_flitdata),                                                  // o:34
  .dst_ready(ir0_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbiea0_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(r1_activity),                                                   // i:1
  .src_req(r1_req),                                                             // i:1
  .src_sop(r1_sop),                                                             // i:1
  .src_eop(r1_eop),                                                             // i:1
  .src_flitdata(r1_flitdata),                                                   // i:24
  .src_ready(r1_ready),                                                         // o:1
  .dst_activity(ir1_activity),                                                  // o:1
  .dst_req(ir1_req),                                                            // o:1
  .dst_sop(ir1_sop),                                                            // o:1
  .dst_eop(ir1_eop),                                                            // o:1
  .dst_flitdata(ir1_flitdata),                                                  // o:24
  .dst_ready(ir1_ready)                                                         // i:1
);
// =======================================================================
// Signal Declarations
// =======================================================================
// Read / Write Address decode hit lines
// logic     $pAddrW int.rawAddr      desc(Read address adjusted to packet address width);
// Sequencer signals
// Read Command header fields
// Read Data + Status signals
// Write Command + Data Signals
// Write status signals
// logic      $pLenW int.rplen;
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbiea0_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
parameter S_HDR = 3'd0;
parameter S_WR = 3'd1;
parameter S_WR_STS = 3'd2;
parameter S_RD_HDR = 3'd3;
parameter S_RD_PLD = 3'd4;
// ============================================
// Clock Gating Logic
// ============================================
assign gclkEn = (int_psel && !int_penable) || if0_req || if1_req || ir0_activity || ir1_activity || ir0_req || ir1_req;
usb4_tc_noc_apbiea0_gcg gcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
assign if0_activity = (int_psel && !int_penable) || (int_psel && int_pwrite);
assign if1_activity = (int_psel && !int_penable) || (int_psel && !int_pwrite);
// =======================================================================
// Decode Read / Write Address and generate hit lines
// =======================================================================
assign rc_rawAddr = int_paddr;
always_comb
begin
  rtmp_did     = 3'd0;
  rtmp_valid   = 1'b0;
  rc_did      = 3'd0;
  rc_sid      = 3'd1;
  rc_mapdAddr = rc_rawAddr;
  if (!int_pwrite && (int_paddr & 32'hC0000) == 32'h0)
    begin
        rtmp_did = 3'd6;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hFFE00) == 32'h40000)
    begin
        rtmp_did = 3'd1;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hF0000) == 32'h50000)
    begin
        rtmp_did = 3'd2;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hF0000) == 32'h60000)
    begin
        rtmp_did = 3'd3;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hF0000) == 32'h70000)
    begin
        rtmp_did = 3'd4;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hFFC00) == 32'h40400)
    begin
        rtmp_did = 3'd5;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
end

assign wcd_rawAddr = int_paddr;
always_comb
begin
  wtmp_did     = 3'd0;
  wtmp_valid   = 1'b0;
  wcd_did      = 3'd0;
  wcd_sid      = 3'd1;
  wcd_mapdAddr = wcd_rawAddr;
  if ( int_pwrite && (int_paddr & 32'hC0000) == 32'h0)
    begin
      wtmp_did = 3'd6;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hFFE00) == 32'h40000)
    begin
      wtmp_did = 3'd1;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hF0000) == 32'h50000)
    begin
      wtmp_did = 3'd2;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hF0000) == 32'h60000)
    begin
      wtmp_did = 3'd3;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hF0000) == 32'h70000)
    begin
      wtmp_did = 3'd4;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hFFC00) == 32'h40400)
    begin
      wtmp_did = 3'd5;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
end

// ============================================
// Target Local Address Translation
// ============================================
// =======================================================================
// Read Command Path Processing
// =======================================================================
// ============================================
// Read Command header field assignments
// ============================================
// ============================================
// Read Command header field packing
// ============================================
assign rpaylen = 3'd4 - (3'(rc_mapdAddr) & 3'd3);
always_comb
begin
  // Set default header to all 0s
  rc_hdr               = {60{1'b0}};
  // Assign over the various fields
  rc_hdr[3:0]    = 4'd4;                                                        // QoS: set to mid qos value
  rc_hdr[6:4]    = rc_did;                                                      // Destination ID
  rc_hdr[7]    = 1'b1;                                                          // SoT: not supporting fragmentation at the moment
  rc_hdr[8]    = 1'b1;                                                          // EoT: not supporting fragmentation at the moment
  rc_hdr[14:9]    = 6'd0;                                                       // Read command
  rc_hdr[17:15]    = rc_sid;                                                    // Initiator ID
  rc_hdr[19:18]    = 2'd0;                                                      // Transaction ID
  rc_hdr[22:20]   = rpaylen;                                                    // Packet length is always one data phase long
  rc_hdr[54:23]   = rc_mapdAddr[31:0];
  rc_hdr[57:55]   = 3'd2;                                                       // Size is log2 of width of bus
  rc_hdr[59:58]  = 2'd1;                                                        // Always incrementing
  // Security attributes
  // User Attributes
end

// =======================================================================
// Write Command and Data Path Processing
// =======================================================================
// ============================================
// Write Command Header field assignments
// ============================================
assign wpaylen = 3'd4 - (3'(wcd_mapdAddr) & 3'd3);
always_comb
begin
  // Set default header to all 0s
  wcd_hdr              = {72{1'b0}};
  // Assign over the various fields
  wcd_hdr[3:0]    = 4'd4;                                                       // QoS: set to mid qos value
  wcd_hdr[6:4]    = wcd_did;                                                    // Destination ID
  wcd_hdr[7]    = 1'b1;                                                         // SoT: not supporting fragmentation at the moment
  wcd_hdr[8]    = 1'b1;                                                         // EoT: not supporting fragmentation at the moment
  wcd_hdr[14:9]    = 6'd2;                                                      // Write command + data
  wcd_hdr[17:15]    = wcd_sid;                                                  // Initiator ID
  wcd_hdr[19:18]    = 2'd0;                                                     // Transaction ID
  wcd_hdr[22:20]   = wpaylen;                                                   // Packet length is always one data phase long
  wcd_hdr[54:23]   = wcd_mapdAddr[31:0];
  wcd_hdr[57:55]   = 3'd2;                                                      // Size is log2 of width of bus
  wcd_hdr[59:58]  = 2'd1;                                                       // Always incrementing
  // Security attributes
  // User Attributes
end

assign wcd_pld = {{int_pstrb[3:0],int_pwdata[31:0]}};
// Write Status Buffer
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      ws_buf[0] <= #1ps 24'd0;
    end
  else
    begin
      if (ws_buf_en[0])
        ws_buf[0] <= #1ps ir1_flitdata;
    end
end

assign ws_buf_en = ws_buf_we << fcnt;
// =======================================================================
// Write Status Path Processing
// =======================================================================
assign ws_bus = {ir1_flitdata };
// ============================================
// Read / Write Command flit sequencer
// ============================================
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    fcnt <= #1ps 1'd0;
  else if (fcnt_en)
    fcnt <= #1ps fcnt_nxt;
end

// Read Data + Status Buffer
// Header Buffer
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rs_buf[0] <= #1ps {34{1'b0}};
      rs_buf[1] <= #1ps {34{1'b0}};
    end
  else
    begin
      if (rs_buf_en[0])
        rs_buf[0] <= #1ps ir0_flitdata;
      if (rs_buf_en[1])
        rs_buf[1] <= #1ps ir0_flitdata;
    end
end

assign rs_buf_en = rs_buf_we << fcnt;
// Create incoming rs.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rs_bus[33:0] = rs_buf[0];
assign rs_bus[67:34] = ((state == S_RD_HDR) && (fcnt == 1'd1)) ? ir0_flitdata : rs_buf[1];
// =======================================================================
// Read Data and Status Path Processing
// =======================================================================
assign rds_bus = {ir0_flitdata };
assign rds_data = {readSeg[31:0]};
assign rds_status = {readSeg[33:32]};
assign readSeg = rds_bus;
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    state <= #1ps S_HDR;
  else
    state <= #1ps state_nxt;
end

// pp: my $condRuW = $ruW;   # Condition read user width - clears effective ruW if NoC packet does not include ruser
always_comb
begin
  fcnt_nxt    = fcnt;
  fcnt_en     = 1'b0;
  state_nxt   = state;
  int_pready  = 1'b0;
  int_prdata  = 32'd0;
  int_pslverr = 1'b0;
  if0_req     = 1'b0;
  if0_sop     = 1'b0;
  if0_eop     = 1'b0;
  if0_flitdata = {36{1'b0}};
  ir1_ready   = 1'b0;
  ws_buf_we   = 1'b0;
  if1_req     = 1'b0;
  if1_sop     = 1'b0;
  if1_eop     = 1'b0;
  if1_flitdata = {60{1'b0}};
  ir0_ready   = 1'b0;
  rs_buf_we  = 1'b0;
  case (state)
    S_HDR:
      begin
        // Slave is being selected for write access
        if (int_psel && int_penable && int_pwrite)
          begin
            if0_req = 1'b1;
            if0_sop = (fcnt == 1'd0);
            // Generate the f0 flit data
            case(fcnt)
              1'd0: if0_flitdata = wcd_hdr[35:0];
              1'd1: if0_flitdata = wcd_hdr[71:36];
              default: if0_flitdata = {36{1'b0}};
            endcase
            // Update the header fragment count and generate the ready back to the ingress pipe stage
            if (int_psel && if0_ready)
              begin
                if (fcnt == 1'd1)
                  begin
                    fcnt_nxt    = 1'd0;
                    fcnt_en     = 1'b1;
                    state_nxt   = S_WR;
                  end
               else
                  begin
                    fcnt_nxt  = fcnt + 1'd1;
                    fcnt_en   = 1'b1;
                   end
              end
          end
        // Slave is being selected for read access
        else if (int_psel && int_penable && !int_pwrite)
          begin
            if1_req     = 1'b1;
            if1_sop     = (fcnt == 1'd0);
            if1_eop     = (fcnt == 1'd0);
            case(fcnt)
              1'd0: if1_flitdata = rc_hdr[59:0];
              default: if1_flitdata = {60{1'b0}};
            endcase
            // Update the header fragment count and generate the ready back to the ingress pipe stage
            // Header transmission is complete
            if (int_psel && if1_ready)
              begin
                if (fcnt == 1'd0)
                  begin
                    fcnt_nxt  = 1'd0;
                    fcnt_en   = 1'b1;
                    state_nxt = S_RD_HDR;
                  end
                // Continuing header transmission
                else
                  begin
                    fcnt_nxt = fcnt + 1'd1;
                    fcnt_en  = 1'b1;
                  end
              end
          end
      end
    S_WR:
      begin
        if0_req = 1'b1;
        if0_eop = (fcnt == 1'd0);
        if0_flitdata = {36{1'b0}};
        if0_flitdata = wcd_pld;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_ready)
          begin
            // Complete data phase is done
            if (fcnt == 1'd0)
              begin
                fcnt_nxt   = 1'd0;
                fcnt_en    = 1'b1;
                state_nxt  = S_WR_STS;
              end
            else
              begin
                fcnt_nxt   = fcnt + 1'd1;
                fcnt_en    = 1'b1;
              end
          end
      end
    S_WR_STS:
      begin
        ir1_ready   = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_req)
          begin
            // Header transmission is complete
            if (fcnt == 1'd0)
              begin
                int_pready  = 1'b1;
                int_pslverr = |ws_bus[23:20];
                fcnt_nxt    = 1'd0;
                fcnt_en     = 1'b1;
                state_nxt   = S_HDR;
              end
            // Continuing header transmission
            else
              begin
                fcnt_nxt  = fcnt + 1'd1;
                fcnt_en   = 1'b1;
                ws_buf_we = 1'b1;
              end
          end
      end
    S_RD_HDR:
      begin
        // Update the header fragment count and generate the ready back to the r0 interface
        ir0_ready = 1'b1;
        if (ir0_req)
          begin
            // Complete read header is done
            if (fcnt == 1'd1)
              begin
                fcnt_nxt   = 1'd0;
                fcnt_en    = 1'b1;
                state_nxt   = S_RD_PLD;
                rs_buf_we = 1'b1;
              end
            else
              begin
                fcnt_nxt   = fcnt + 1'd1;
                fcnt_en    = 1'b1;
                rs_buf_we = 1'b1;
              end
          end
      end
    S_RD_PLD:
      begin
        // Update the header fragment count and generate the ready back to the r0 interface
        ir0_ready = 1'b1;
        if (ir0_req)
          begin
            // Complete read header is done
            if (fcnt == 1'd0)
              begin
                int_pready  = 1'b1;
                int_pslverr = |rds_status;
                int_prdata  = rds_data;
                fcnt_nxt    = 1'd0;
                fcnt_en     = 1'b1;
                state_nxt   = S_HDR;
              end
            else
              begin
                fcnt_nxt   = fcnt + 1'd1;
                fcnt_en    = 1'b1;
              end
          end
      end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_ipipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire     [31:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  output logic           src_pslverr,                                           // Slave error
  // dst
  output logic    [31:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata,                                            // Read data
  input  wire            dst_pslverr                                            // Slave error
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbiea0_ipipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
assign src_pslverr = dst_pslverr;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_ipipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea0_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea0_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea0_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea0_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea0_gcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1 (
  input  wire            clk,
  input  wire            rst_n,
  // s
  input  wire     [31:0] s_paddr,                                               // Address
  input  wire            s_psel,                                                // Select
  input  wire            s_penable,                                             // Enable
  input  wire            s_pwrite,                                              // Write not read
  input  wire     [31:0] s_pwdata,                                              // Write data
  input  wire      [3:0] s_pstrb,                                               // Write strobes
  output logic           s_pready,                                              // Ready
  output logic    [31:0] s_prdata,                                              // Read data
  output logic           s_pslverr,                                             // Slave error
  // f0
  output logic           f0_activity,                                           // Upcoming activity indicator
  output logic           f0_req,                                                // Flit transfer request
  output logic           f0_sop,                                                // Start of packet indicator
  output logic           f0_eop,                                                // End of packet indicator
  output logic    [35:0] f0_flitdata,                                           // Flit data
  input  wire            f0_ready,                                              // Flit transfer ready
  // f1
  output logic           f1_activity,                                           // Upcoming activity indicator
  output logic           f1_req,                                                // Flit transfer request
  output logic           f1_sop,                                                // Start of packet indicator
  output logic           f1_eop,                                                // End of packet indicator
  output logic    [59:0] f1_flitdata,                                           // Flit data
  input  wire            f1_ready,                                              // Flit transfer ready
  // r0
  input  wire            r0_activity,                                           // Upcoming activity indicator
  input  wire            r0_req,                                                // Flit transfer request
  input  wire            r0_sop,                                                // Start of packet indicator
  input  wire            r0_eop,                                                // End of packet indicator
  input  wire     [33:0] r0_flitdata,                                           // Flit data
  output logic           r0_ready,                                              // Flit transfer ready
  // r1
  input  wire            r1_activity,                                           // Upcoming activity indicator
  input  wire            r1_req,                                                // Flit transfer request
  input  wire            r1_sop,                                                // Start of packet indicator
  input  wire            r1_eop,                                                // End of packet indicator
  input  wire     [23:0] r1_flitdata,                                           // Flit data
  output logic           r1_ready                                               // Flit transfer ready
);

logic    [31:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           int_pslverr;                                                    // Slave error
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic     [2:0] rc_did;
logic     [2:0] rc_sid;
logic    [59:0] rc_hdr;
logic    [31:0] rc_rawAddr;
logic    [31:0] rc_mapdAddr;
logic           rs_buf_we;
logic    [67:0] rs_bus;
logic    [33:0] rds_bus;
logic    [31:0] rds_data;
logic     [1:0] rds_status;
logic     [2:0] wcd_did;
logic     [2:0] wcd_sid;
logic    [71:0] wcd_hdr;
logic    [35:0] wcd_pld;
logic    [31:0] wcd_rawAddr;
logic    [31:0] wcd_mapdAddr;
logic           ws_buf_we;
logic    [23:0] ws_bus;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           gclk;
logic           gclkAct;
logic           gclkEn;
logic     [2:0] rtmp_did;
logic           rtmp_valid;
logic     [2:0] wtmp_did;
logic           wtmp_valid;
logic     [2:0] rpaylen;
logic     [2:0] wpaylen;
logic    [23:0] ws_buf [0:0];
logic     [0:0] ws_buf_en;
logic     [0:0] fcnt;
logic     [0:0] fcnt_nxt;
logic     [0:0] fcnt_en;
logic    [33:0] rs_buf [1:0];
logic     [1:0] rs_buf_en;
logic    [33:0] readSeg;
logic     [2:0] state;
logic     [2:0] state_nxt;
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Initiator Ports (APB subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Ingress APB Pipeline Component
usb4_tc_noc_apbiea1_ipipe ipipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(s_paddr),                                                          // i:32
  .src_psel(s_psel),                                                            // i:1
  .src_penable(s_penable),                                                      // i:1
  .src_pwrite(s_pwrite),                                                        // i:1
  .src_pwdata(s_pwdata),                                                        // i:32
  .src_pstrb(s_pstrb),                                                          // i:4
  .src_pready(s_pready),                                                        // o:1
  .src_prdata(s_prdata),                                                        // o:32
  .src_pslverr(s_pslverr),                                                      // o:1
  .dst_paddr(int_paddr),                                                        // o:32
  .dst_psel(int_psel),                                                          // o:1
  .dst_penable(int_penable),                                                    // o:1
  .dst_pwrite(int_pwrite),                                                      // o:1
  .dst_pwdata(int_pwdata),                                                      // o:32
  .dst_pstrb(int_pstrb),                                                        // o:4
  .dst_pready(int_pready),                                                      // i:1
  .dst_prdata(int_prdata),                                                      // i:32
  .dst_pslverr(int_pslverr)                                                     // i:1
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbiea1_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(if0_activity),                                                  // i:1
  .src_req(if0_req),                                                            // i:1
  .src_sop(if0_sop),                                                            // i:1
  .src_eop(if0_eop),                                                            // i:1
  .src_flitdata(if0_flitdata),                                                  // i:36
  .src_ready(if0_ready),                                                        // o:1
  .dst_activity(f0_activity),                                                   // o:1
  .dst_req(f0_req),                                                             // o:1
  .dst_sop(f0_sop),                                                             // o:1
  .dst_eop(f0_eop),                                                             // o:1
  .dst_flitdata(f0_flitdata),                                                   // o:36
  .dst_ready(f0_ready)                                                          // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbiea1_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(if1_activity),                                                  // i:1
  .src_req(if1_req),                                                            // i:1
  .src_sop(if1_sop),                                                            // i:1
  .src_eop(if1_eop),                                                            // i:1
  .src_flitdata(if1_flitdata),                                                  // i:60
  .src_ready(if1_ready),                                                        // o:1
  .dst_activity(f1_activity),                                                   // o:1
  .dst_req(f1_req),                                                             // o:1
  .dst_sop(f1_sop),                                                             // o:1
  .dst_eop(f1_eop),                                                             // o:1
  .dst_flitdata(f1_flitdata),                                                   // o:60
  .dst_ready(f1_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbiea1_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(r0_activity),                                                   // i:1
  .src_req(r0_req),                                                             // i:1
  .src_sop(r0_sop),                                                             // i:1
  .src_eop(r0_eop),                                                             // i:1
  .src_flitdata(r0_flitdata),                                                   // i:34
  .src_ready(r0_ready),                                                         // o:1
  .dst_activity(ir0_activity),                                                  // o:1
  .dst_req(ir0_req),                                                            // o:1
  .dst_sop(ir0_sop),                                                            // o:1
  .dst_eop(ir0_eop),                                                            // o:1
  .dst_flitdata(ir0_flitdata),                                                  // o:34
  .dst_ready(ir0_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbiea1_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(r1_activity),                                                   // i:1
  .src_req(r1_req),                                                             // i:1
  .src_sop(r1_sop),                                                             // i:1
  .src_eop(r1_eop),                                                             // i:1
  .src_flitdata(r1_flitdata),                                                   // i:24
  .src_ready(r1_ready),                                                         // o:1
  .dst_activity(ir1_activity),                                                  // o:1
  .dst_req(ir1_req),                                                            // o:1
  .dst_sop(ir1_sop),                                                            // o:1
  .dst_eop(ir1_eop),                                                            // o:1
  .dst_flitdata(ir1_flitdata),                                                  // o:24
  .dst_ready(ir1_ready)                                                         // i:1
);
// =======================================================================
// Signal Declarations
// =======================================================================
// Read / Write Address decode hit lines
// logic     $pAddrW int.rawAddr      desc(Read address adjusted to packet address width);
// Sequencer signals
// Read Command header fields
// Read Data + Status signals
// Write Command + Data Signals
// Write status signals
// logic      $pLenW int.rplen;
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbiea1_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
parameter S_HDR = 3'd0;
parameter S_WR = 3'd1;
parameter S_WR_STS = 3'd2;
parameter S_RD_HDR = 3'd3;
parameter S_RD_PLD = 3'd4;
// ============================================
// Clock Gating Logic
// ============================================
assign gclkEn = (int_psel && !int_penable) || if0_req || if1_req || ir0_activity || ir1_activity || ir0_req || ir1_req;
usb4_tc_noc_apbiea1_gcg gcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
assign if0_activity = (int_psel && !int_penable) || (int_psel && int_pwrite);
assign if1_activity = (int_psel && !int_penable) || (int_psel && !int_pwrite);
// =======================================================================
// Decode Read / Write Address and generate hit lines
// =======================================================================
assign rc_rawAddr = int_paddr;
always_comb
begin
  rtmp_did     = 3'd0;
  rtmp_valid   = 1'b0;
  rc_did      = 3'd0;
  rc_sid      = 3'd2;
  rc_mapdAddr = rc_rawAddr;
  if (!int_pwrite && (int_paddr & 32'hC0000) == 32'h0)
    begin
        rtmp_did = 3'd6;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hFFE00) == 32'h40000)
    begin
        rtmp_did = 3'd1;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hF0000) == 32'h50000)
    begin
        rtmp_did = 3'd2;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hF0000) == 32'h60000)
    begin
        rtmp_did = 3'd3;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hF0000) == 32'h70000)
    begin
        rtmp_did = 3'd4;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hFFC00) == 32'h40400)
    begin
        rtmp_did = 3'd5;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
  if (!int_pwrite && (int_paddr & 32'hFF000) == 32'h80000)
    begin
        rtmp_did = 3'd0;
        rtmp_valid = 1'b0;
        rtmp_valid = 1'b1;
        if( rtmp_valid )
          begin
            rc_did = rtmp_did;
          end
        else
          begin
            rc_did      = 3'd0;
          end
      rc_mapdAddr = rc_rawAddr;
    end
end

assign wcd_rawAddr = int_paddr;
always_comb
begin
  wtmp_did     = 3'd0;
  wtmp_valid   = 1'b0;
  wcd_did      = 3'd0;
  wcd_sid      = 3'd2;
  wcd_mapdAddr = wcd_rawAddr;
  if ( int_pwrite && (int_paddr & 32'hC0000) == 32'h0)
    begin
      wtmp_did = 3'd6;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hFFE00) == 32'h40000)
    begin
      wtmp_did = 3'd1;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hF0000) == 32'h50000)
    begin
      wtmp_did = 3'd2;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hF0000) == 32'h60000)
    begin
      wtmp_did = 3'd3;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hF0000) == 32'h70000)
    begin
      wtmp_did = 3'd4;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hFFC00) == 32'h40400)
    begin
      wtmp_did = 3'd5;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
  if ( int_pwrite && (int_paddr & 32'hFF000) == 32'h80000)
    begin
      wtmp_did = 3'd0;
      wtmp_valid = 1'b0;
      wtmp_valid = 1'b1;
      if( wtmp_valid )
        begin
          wcd_did = wtmp_did;
        end
      else
        begin
          wcd_did      = 3'd0;
        end
      wcd_mapdAddr = wcd_rawAddr;
    end
end

// ============================================
// Target Local Address Translation
// ============================================
// =======================================================================
// Read Command Path Processing
// =======================================================================
// ============================================
// Read Command header field assignments
// ============================================
// ============================================
// Read Command header field packing
// ============================================
assign rpaylen = 3'd4 - (3'(rc_mapdAddr) & 3'd3);
always_comb
begin
  // Set default header to all 0s
  rc_hdr               = {60{1'b0}};
  // Assign over the various fields
  rc_hdr[3:0]    = 4'd4;                                                        // QoS: set to mid qos value
  rc_hdr[6:4]    = rc_did;                                                      // Destination ID
  rc_hdr[7]    = 1'b1;                                                          // SoT: not supporting fragmentation at the moment
  rc_hdr[8]    = 1'b1;                                                          // EoT: not supporting fragmentation at the moment
  rc_hdr[14:9]    = 6'd0;                                                       // Read command
  rc_hdr[17:15]    = rc_sid;                                                    // Initiator ID
  rc_hdr[19:18]    = 2'd0;                                                      // Transaction ID
  rc_hdr[22:20]   = rpaylen;                                                    // Packet length is always one data phase long
  rc_hdr[54:23]   = rc_mapdAddr[31:0];
  rc_hdr[57:55]   = 3'd2;                                                       // Size is log2 of width of bus
  rc_hdr[59:58]  = 2'd1;                                                        // Always incrementing
  // Security attributes
  // User Attributes
end

// =======================================================================
// Write Command and Data Path Processing
// =======================================================================
// ============================================
// Write Command Header field assignments
// ============================================
assign wpaylen = 3'd4 - (3'(wcd_mapdAddr) & 3'd3);
always_comb
begin
  // Set default header to all 0s
  wcd_hdr              = {72{1'b0}};
  // Assign over the various fields
  wcd_hdr[3:0]    = 4'd4;                                                       // QoS: set to mid qos value
  wcd_hdr[6:4]    = wcd_did;                                                    // Destination ID
  wcd_hdr[7]    = 1'b1;                                                         // SoT: not supporting fragmentation at the moment
  wcd_hdr[8]    = 1'b1;                                                         // EoT: not supporting fragmentation at the moment
  wcd_hdr[14:9]    = 6'd2;                                                      // Write command + data
  wcd_hdr[17:15]    = wcd_sid;                                                  // Initiator ID
  wcd_hdr[19:18]    = 2'd0;                                                     // Transaction ID
  wcd_hdr[22:20]   = wpaylen;                                                   // Packet length is always one data phase long
  wcd_hdr[54:23]   = wcd_mapdAddr[31:0];
  wcd_hdr[57:55]   = 3'd2;                                                      // Size is log2 of width of bus
  wcd_hdr[59:58]  = 2'd1;                                                       // Always incrementing
  // Security attributes
  // User Attributes
end

assign wcd_pld = {{int_pstrb[3:0],int_pwdata[31:0]}};
// Write Status Buffer
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      ws_buf[0] <= #1ps 24'd0;
    end
  else
    begin
      if (ws_buf_en[0])
        ws_buf[0] <= #1ps ir1_flitdata;
    end
end

assign ws_buf_en = ws_buf_we << fcnt;
// =======================================================================
// Write Status Path Processing
// =======================================================================
assign ws_bus = {ir1_flitdata };
// ============================================
// Read / Write Command flit sequencer
// ============================================
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    fcnt <= #1ps 1'd0;
  else if (fcnt_en)
    fcnt <= #1ps fcnt_nxt;
end

// Read Data + Status Buffer
// Header Buffer
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rs_buf[0] <= #1ps {34{1'b0}};
      rs_buf[1] <= #1ps {34{1'b0}};
    end
  else
    begin
      if (rs_buf_en[0])
        rs_buf[0] <= #1ps ir0_flitdata;
      if (rs_buf_en[1])
        rs_buf[1] <= #1ps ir0_flitdata;
    end
end

assign rs_buf_en = rs_buf_we << fcnt;
// Create incoming rs.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rs_bus[33:0] = rs_buf[0];
assign rs_bus[67:34] = ((state == S_RD_HDR) && (fcnt == 1'd1)) ? ir0_flitdata : rs_buf[1];
// =======================================================================
// Read Data and Status Path Processing
// =======================================================================
assign rds_bus = {ir0_flitdata };
assign rds_data = {readSeg[31:0]};
assign rds_status = {readSeg[33:32]};
assign readSeg = rds_bus;
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    state <= #1ps S_HDR;
  else
    state <= #1ps state_nxt;
end

// pp: my $condRuW = $ruW;   # Condition read user width - clears effective ruW if NoC packet does not include ruser
always_comb
begin
  fcnt_nxt    = fcnt;
  fcnt_en     = 1'b0;
  state_nxt   = state;
  int_pready  = 1'b0;
  int_prdata  = 32'd0;
  int_pslverr = 1'b0;
  if0_req     = 1'b0;
  if0_sop     = 1'b0;
  if0_eop     = 1'b0;
  if0_flitdata = {36{1'b0}};
  ir1_ready   = 1'b0;
  ws_buf_we   = 1'b0;
  if1_req     = 1'b0;
  if1_sop     = 1'b0;
  if1_eop     = 1'b0;
  if1_flitdata = {60{1'b0}};
  ir0_ready   = 1'b0;
  rs_buf_we  = 1'b0;
  case (state)
    S_HDR:
      begin
        // Slave is being selected for write access
        if (int_psel && int_penable && int_pwrite)
          begin
            if0_req = 1'b1;
            if0_sop = (fcnt == 1'd0);
            // Generate the f0 flit data
            case(fcnt)
              1'd0: if0_flitdata = wcd_hdr[35:0];
              1'd1: if0_flitdata = wcd_hdr[71:36];
              default: if0_flitdata = {36{1'b0}};
            endcase
            // Update the header fragment count and generate the ready back to the ingress pipe stage
            if (int_psel && if0_ready)
              begin
                if (fcnt == 1'd1)
                  begin
                    fcnt_nxt    = 1'd0;
                    fcnt_en     = 1'b1;
                    state_nxt   = S_WR;
                  end
               else
                  begin
                    fcnt_nxt  = fcnt + 1'd1;
                    fcnt_en   = 1'b1;
                   end
              end
          end
        // Slave is being selected for read access
        else if (int_psel && int_penable && !int_pwrite)
          begin
            if1_req     = 1'b1;
            if1_sop     = (fcnt == 1'd0);
            if1_eop     = (fcnt == 1'd0);
            case(fcnt)
              1'd0: if1_flitdata = rc_hdr[59:0];
              default: if1_flitdata = {60{1'b0}};
            endcase
            // Update the header fragment count and generate the ready back to the ingress pipe stage
            // Header transmission is complete
            if (int_psel && if1_ready)
              begin
                if (fcnt == 1'd0)
                  begin
                    fcnt_nxt  = 1'd0;
                    fcnt_en   = 1'b1;
                    state_nxt = S_RD_HDR;
                  end
                // Continuing header transmission
                else
                  begin
                    fcnt_nxt = fcnt + 1'd1;
                    fcnt_en  = 1'b1;
                  end
              end
          end
      end
    S_WR:
      begin
        if0_req = 1'b1;
        if0_eop = (fcnt == 1'd0);
        if0_flitdata = {36{1'b0}};
        if0_flitdata = wcd_pld;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_ready)
          begin
            // Complete data phase is done
            if (fcnt == 1'd0)
              begin
                fcnt_nxt   = 1'd0;
                fcnt_en    = 1'b1;
                state_nxt  = S_WR_STS;
              end
            else
              begin
                fcnt_nxt   = fcnt + 1'd1;
                fcnt_en    = 1'b1;
              end
          end
      end
    S_WR_STS:
      begin
        ir1_ready   = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_req)
          begin
            // Header transmission is complete
            if (fcnt == 1'd0)
              begin
                int_pready  = 1'b1;
                int_pslverr = |ws_bus[23:20];
                fcnt_nxt    = 1'd0;
                fcnt_en     = 1'b1;
                state_nxt   = S_HDR;
              end
            // Continuing header transmission
            else
              begin
                fcnt_nxt  = fcnt + 1'd1;
                fcnt_en   = 1'b1;
                ws_buf_we = 1'b1;
              end
          end
      end
    S_RD_HDR:
      begin
        // Update the header fragment count and generate the ready back to the r0 interface
        ir0_ready = 1'b1;
        if (ir0_req)
          begin
            // Complete read header is done
            if (fcnt == 1'd1)
              begin
                fcnt_nxt   = 1'd0;
                fcnt_en    = 1'b1;
                state_nxt   = S_RD_PLD;
                rs_buf_we = 1'b1;
              end
            else
              begin
                fcnt_nxt   = fcnt + 1'd1;
                fcnt_en    = 1'b1;
                rs_buf_we = 1'b1;
              end
          end
      end
    S_RD_PLD:
      begin
        // Update the header fragment count and generate the ready back to the r0 interface
        ir0_ready = 1'b1;
        if (ir0_req)
          begin
            // Complete read header is done
            if (fcnt == 1'd0)
              begin
                int_pready  = 1'b1;
                int_pslverr = |rds_status;
                int_prdata  = rds_data;
                fcnt_nxt    = 1'd0;
                fcnt_en     = 1'b1;
                state_nxt   = S_HDR;
              end
            else
              begin
                fcnt_nxt   = fcnt + 1'd1;
                fcnt_en    = 1'b1;
              end
          end
      end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_ipipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire     [31:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  output logic           src_pslverr,                                           // Slave error
  // dst
  output logic    [31:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata,                                            // Read data
  input  wire            dst_pslverr                                            // Slave error
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbiea1_ipipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
assign src_pslverr = dst_pslverr;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_ipipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea1_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea1_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea1_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbiea1_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbiea1_gcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0 (
  input  wire            clk,
  input  wire            rst_n,
  // t
  output logic     [8:0] t_paddr,                                               // Address
  output logic           t_psel,                                                // Select
  output logic           t_penable,                                             // Enable
  output logic           t_pwrite,                                              // Write not read
  output logic    [31:0] t_pwdata,                                              // Write data
  output logic     [3:0] t_pstrb,                                               // Write strobes
  input  wire            t_pready,                                              // Ready
  input  wire     [31:0] t_prdata,                                              // Read data
  // f0
  input  wire            f0_activity,                                           // Upcoming activity indicator
  input  wire            f0_req,                                                // Flit transfer request
  input  wire            f0_sop,                                                // Start of packet indicator
  input  wire            f0_eop,                                                // End of packet indicator
  input  wire     [35:0] f0_flitdata,                                           // Flit data
  output logic           f0_ready,                                              // Flit transfer ready
  // f1
  input  wire            f1_activity,                                           // Upcoming activity indicator
  input  wire            f1_req,                                                // Flit transfer request
  input  wire            f1_sop,                                                // Start of packet indicator
  input  wire            f1_eop,                                                // End of packet indicator
  input  wire     [59:0] f1_flitdata,                                           // Flit data
  output logic           f1_ready,                                              // Flit transfer ready
  // r0
  output logic           r0_activity,                                           // Upcoming activity indicator
  output logic           r0_req,                                                // Flit transfer request
  output logic           r0_sop,                                                // Start of packet indicator
  output logic           r0_eop,                                                // End of packet indicator
  output logic    [33:0] r0_flitdata,                                           // Flit data
  input  wire            r0_ready,                                              // Flit transfer ready
  // r1
  output logic           r1_activity,                                           // Upcoming activity indicator
  output logic           r1_req,                                                // Flit transfer request
  output logic           r1_sop,                                                // Start of packet indicator
  output logic           r1_eop,                                                // End of packet indicator
  output logic    [23:0] r1_flitdata,                                           // Flit data
  input  wire            r1_ready                                               // Flit transfer ready
);

logic     [8:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic           wr_req;
logic           wr_ready;
logic           wr_last;
logic    [31:0] wr_data;
logic     [3:0] wr_strb;
logic           wc_buf_we;
logic    [71:0] wc_bus;
logic     [2:0] wc_sid;
logic     [2:0] wc_did;
logic     [1:0] wc_id;
logic    [31:0] wc_addr;
logic     [7:0] wc_len;
logic     [2:0] wc_rawsize;
logic     [2:0] wc_size;
logic     [1:0] wc_burst;
logic     [3:0] wc_qos;
logic     [2:0] wc_plen;
logic     [2:0] wc_prot;
logic           wcd_transinfo_en;
logic           wcd_transinfo_rdy;
logic           wf_req;
logic           wf_eop;
logic    [35:0] wf_flitdata;
logic           wf_ready;
logic    [23:0] ws_hdr;
logic           int_awvalid;
logic    [67:0] rds_hdr;
logic           rd_req;
logic           rd_ready;
logic           rd_last;
logic           rc_buf_we;
logic    [59:0] rc_bus;
logic     [2:0] rc_sid;
logic     [2:0] rc_did;
logic     [1:0] rc_id;
logic    [31:0] rc_addr;
logic     [2:0] rc_rawsize;
logic     [2:0] rc_size;
logic     [1:0] rc_burst;
logic     [3:0] rc_qos;
logic     [2:0] rc_plen;
logic     [2:0] rc_prot;
logic           rf_req;
logic           rf_eop;
logic    [33:0] rf_flitdata;
logic           rf_ready;
logic           rds_transinfo_we;
logic           rds_transinfo_rdy;
logic           int_arvalid;
logic    [11:0] wc_addr_unpack;
logic    [11:0] rc_addr_pack;
logic     [2:0] int_pprot;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           apbclk;
logic           apbclkAct;
logic           int_apbactivity;
logic           wcclk;
logic           wcclkAct;
wire            int_awactivity;
logic           wdclk;
logic           wdclkAct;
logic           int_wactivity;
logic           rcclk;
logic           rcclkAct;
logic           int_aractivity;
logic           rdclk;
logic           rdclkAct;
logic           rdclkEn;
logic           wrDone;
logic     [0:0] wr_cnt;
logic     [0:0] wr_cnt_nxt;
logic     [0:0] wr_cnt_en;
logic     [1:0] wr_state;
logic     [1:0] wr_state_nxt;
logic     [0:0] wr_state_en;
logic    [35:0] wc_buf [1:0];
logic     [1:0] wc_buf_en;
logic           int_pslverr;
logic     [0:0] rc_cnt;
logic     [0:0] rc_cnt_nxt;
logic     [0:0] rc_cnt_en;
logic           pslverr_w;
logic    [31:0] prdata;
logic     [1:0] rd_state;
logic     [1:0] rd_state_nxt;
logic     [0:0] rd_state_en;
logic    [59:0] rc_buf [0:0];
logic     [0:0] rc_buf_en;
logic           Narrow_Req;
logic     [1:0] apb_state;
logic     [1:0] apb_state_nxt;
logic     [0:0] apb_state_en;
logic     [0:0] apb_wrarb;
logic     [0:0] apb_wrarb_nxt;
logic     [0:0] apb_wrarb_en;
// ========================================================================//
// Parameter Declarations
// ========================================================================//
// ========================================================================//
// Process parameters and create local derived variables
// ========================================================================//
// ========================================================================//
// Define module I/O
// ========================================================================//
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Target Interface(s) (APB manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Egress APB Pipeline Component
usb4_tc_noc_apbtea0_epipe epipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(int_paddr),                                                        // i:9
  .src_psel(int_psel),                                                          // i:1
  .src_penable(int_penable),                                                    // i:1
  .src_pwrite(int_pwrite),                                                      // i:1
  .src_pwdata(int_pwdata),                                                      // i:32
  .src_pstrb(int_pstrb),                                                        // i:4
  .src_pready(int_pready),                                                      // o:1
  .src_prdata(int_prdata),                                                      // o:32
  .dst_paddr(t_paddr),                                                          // o:9
  .dst_psel(t_psel),                                                            // o:1
  .dst_penable(t_penable),                                                      // o:1
  .dst_pwrite(t_pwrite),                                                        // o:1
  .dst_pwdata(t_pwdata),                                                        // o:32
  .dst_pstrb(t_pstrb),                                                          // o:4
  .dst_pready(t_pready),                                                        // i:1
  .dst_prdata(t_prdata)                                                         // i:32
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea0_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f0_activity),                                                   // i:1
  .src_req(f0_req),                                                             // i:1
  .src_sop(f0_sop),                                                             // i:1
  .src_eop(f0_eop),                                                             // i:1
  .src_flitdata(f0_flitdata),                                                   // i:36
  .src_ready(f0_ready),                                                         // o:1
  .dst_activity(if0_activity),                                                  // o:1
  .dst_req(if0_req),                                                            // o:1
  .dst_sop(if0_sop),                                                            // o:1
  .dst_eop(if0_eop),                                                            // o:1
  .dst_flitdata(if0_flitdata),                                                  // o:36
  .dst_ready(if0_ready)                                                         // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea0_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f1_activity),                                                   // i:1
  .src_req(f1_req),                                                             // i:1
  .src_sop(f1_sop),                                                             // i:1
  .src_eop(f1_eop),                                                             // i:1
  .src_flitdata(f1_flitdata),                                                   // i:60
  .src_ready(f1_ready),                                                         // o:1
  .dst_activity(if1_activity),                                                  // o:1
  .dst_req(if1_req),                                                            // o:1
  .dst_sop(if1_sop),                                                            // o:1
  .dst_eop(if1_eop),                                                            // o:1
  .dst_flitdata(if1_flitdata),                                                  // o:60
  .dst_ready(if1_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea0_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir0_activity),                                                  // i:1
  .src_req(ir0_req),                                                            // i:1
  .src_sop(ir0_sop),                                                            // i:1
  .src_eop(ir0_eop),                                                            // i:1
  .src_flitdata(ir0_flitdata),                                                  // i:34
  .src_ready(ir0_ready),                                                        // o:1
  .dst_activity(r0_activity),                                                   // o:1
  .dst_req(r0_req),                                                             // o:1
  .dst_sop(r0_sop),                                                             // o:1
  .dst_eop(r0_eop),                                                             // o:1
  .dst_flitdata(r0_flitdata),                                                   // o:34
  .dst_ready(r0_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea0_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir1_activity),                                                  // i:1
  .src_req(ir1_req),                                                            // i:1
  .src_sop(ir1_sop),                                                            // i:1
  .src_eop(ir1_eop),                                                            // i:1
  .src_flitdata(ir1_flitdata),                                                  // i:24
  .src_ready(ir1_ready),                                                        // o:1
  .dst_activity(r1_activity),                                                   // o:1
  .dst_req(r1_req),                                                             // o:1
  .dst_sop(r1_sop),                                                             // o:1
  .dst_eop(r1_eop),                                                             // o:1
  .dst_flitdata(r1_flitdata),                                                   // o:24
  .dst_ready(r1_ready)                                                          // i:1
);
// =======================================================================
// Signal declarations
// =======================================================================
// Write Command + Data Sequencer Signals
// Write Command Signals
// Write Response Fields
// Read Data + Status fields
// Read Data + Status Flit Sequencer Signals
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea0_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign int_apbactivity = int_awactivity || int_aractivity;
usb4_tc_noc_apbtea0_apbcg apbcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_apbactivity),                                                      // i:1
  .clkOut(apbclk),                                                              // o:1
  .isActive(apbclkAct)                                                          // o:1
);
assign int_awactivity = if0_activity || if0_req || int_awvalid || ir1_req || wr_req;
usb4_tc_noc_apbtea0_wccg wccg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_awactivity),                                                       // i:1
  .clkOut(wcclk),                                                               // o:1
  .isActive(wcclkAct)                                                           // o:1
);
assign int_wactivity = if0_activity || if0_req || !wcd_transinfo_rdy || int_awvalid;
usb4_tc_noc_apbtea0_wdcg wdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_wactivity),                                                        // i:1
  .clkOut(wdclk),                                                               // o:1
  .isActive(wdclkAct)                                                           // o:1
);
assign ir1_activity = ir1_req;
assign int_aractivity = if1_activity || if1_req || ir0_req || rd_req;
usb4_tc_noc_apbtea0_f1cg f1cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_aractivity),                                                       // i:1
  .clkOut(rcclk),                                                               // o:1
  .isActive(rcclkAct)                                                           // o:1
);
assign ir0_activity = ir0_req;
assign rdclkEn = ir0_activity || if1_activity || if1_req || !rds_transinfo_rdy;
usb4_tc_noc_apbtea0_rdcg rdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(rdclkEn),                                                              // i:1
  .clkOut(rdclk),                                                               // o:1
  .isActive(rdclkAct)                                                           // o:1
);
// =======================================================================
// Write Processing
// =======================================================================
assign wrDone = wr_last && int_penable && int_pwrite && int_pready;
parameter S_WR_HDR = 2'd0;
parameter S_WR_DATA = 2'd1;
parameter S_WR_WAIT = 2'd2;
parameter S_WR_STS = 2'd3;
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign wc_bus[35:0] = wc_buf[0];
assign wc_bus[71:36] = ((wr_state == 2'b00) && (wr_cnt >= 1'd1)) ? if0_flitdata : wc_buf[1];
// Current Flit Count
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_cnt <= #1ps 1'd0;
  else if (wr_cnt_en)
    wr_cnt <= #1ps wr_cnt_nxt;
end

// Write State Machine State
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_state <= #1ps S_WR_HDR;
  else if (wr_state_en)
    wr_state <= #1ps wr_state_nxt;
end

// Write Command Packing Buffer
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      wc_buf[0] <= #1ps {36{1'b0}};
      wc_buf[1] <= #1ps {36{1'b0}};
    end
  else
    begin
      if (wc_buf_en[0])
        wc_buf[0] <= #1ps if0_flitdata;
      if (wc_buf_en[1])
        wc_buf[1] <= #1ps if0_flitdata;
    end
end

assign wc_buf_en = wc_buf_we << wr_cnt;
always_comb
begin
  // Defaults
  if0_ready    = 1'b0;
  ir1_req      = 1'b0;
  ir1_sop      = 1'b0;
  ir1_eop      = 1'b0;
  ir1_flitdata = {24{1'b0}};
  wr_cnt_nxt   = wr_cnt;
  wr_state_nxt = wr_state;
  wcd_transinfo_en = 1'b0;
  wf_req       = 1'b0;
  wf_eop       = 1'b0;
  wf_flitdata  = {36{1'b0}};
  // Write enables
  wc_buf_we    = 1'b0;
  wr_cnt_en    = 1'b0;
  wr_state_en  = 1'b0;
  int_awvalid   = 1'b0;
  case (wr_state)
    S_WR_HDR:
      begin
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_req)
          begin
            if0_ready    = 1'b1;
            // Header transmission is complete
            if (wr_cnt == 1'd1)
              begin
                int_awvalid = wcd_transinfo_rdy;
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wc_buf_we    = 1'b1;
                wcd_transinfo_en = 1'b1;
                wr_state_nxt = S_WR_DATA;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
                wc_buf_we  = 1'b1;
              end
          end
      end
   S_WR_DATA:
      begin
        wf_req      = if0_req;
        wf_eop      = if0_eop;
        wf_flitdata = if0_flitdata;
        if0_ready   = wf_ready;
        if (if0_req && wf_ready && if0_eop)
          begin
            wr_state_nxt = S_WR_WAIT;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_WAIT:
      begin
        if (wr_req && wr_ready && wr_last)
          begin
            wr_state_nxt = S_WR_STS;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_STS:
      begin
        ir1_req   = 1'b1;
        ir1_sop   = (wr_cnt == 1'd0);
        ir1_eop   = (wr_cnt == 1'd0);
        case(wr_cnt)
          1'd0: ir1_flitdata = ws_hdr[23:0];
          default: ir1_flitdata = {24{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_ready)
          begin
            // Header transmission is complete
            if (wr_cnt == 1'd0)
              begin
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wr_state_nxt = S_WR_HDR;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
              end
          end
      end
  endcase
end

 always_ff @(posedge wcclk) assert ( (frst_n===1'b0) || (int_awvalid == 1'b0) || (wc_burst != 2'b00) || ( {{(32-3){1'b0}},wc_plen} <= (32<<1) )) else $error("ERROR usb4_tc_noc_apbtea0 : %0t : Write data burst request is larger than TEA can handle. Write data burst size(wplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,wc_plen,(32<<1) );
usb4_tc_noc_apbtea0_wdunpack wdunpack (
  .clk(wdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .wtr_req(wcd_transinfo_en),                                                   // i:1
  .wtr_rdy(wcd_transinfo_rdy),                                                  // o:1
  .wtr_size(wc_size),                                                           // i:3
  .wtr_burst(wc_burst),                                                         // i:2
  .wtr_addrlsb(wc_addr[11:0]),                                                  // i:12
  .wtr_plen(wc_plen),                                                           // i:3
  .w_valid(wr_req),                                                             // o:1
  .w_data(wr_data),                                                             // o:32
  .w_strb(wr_strb),                                                             // o:4
  .w_last(wr_last),                                                             // o:1
  .w_ready(wr_ready),                                                           // i:1
  .f_req(wf_req),                                                               // i:1
  .f_eop(wf_eop),                                                               // i:1
  .f_flitdata(wf_flitdata),                                                     // i:36
  .f_ready(wf_ready),                                                           // o:1
  .wtr_addrlsb_out(wc_addr_unpack)                                              // o:12
);
// Write Command + Data Signal Unpacking
assign wc_sid = wc_bus[17:15];
assign wc_did = wc_bus[6:4];
assign wc_id = wc_bus[19:18];
assign wc_addr = wc_bus[54:23];
assign wc_qos = wc_bus[3:0];
assign wc_plen = wc_bus[22:20];
assign wc_prot = 3'd0;
assign wc_rawsize = wc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign wc_size = (wc_rawsize > 3'd2) ? 3'd2 : wc_rawsize;
assign wc_burst = wc_bus[59:58];
// =======================================================================
// Write Response Path Processing
// =======================================================================
// ============================================
// Write Response header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  ws_hdr            = {24{1'b0}};
  // Assign over the various fields
  ws_hdr[3:0]  = wc_qos;                                                        // loopback QoS from write command
  ws_hdr[6:4]  = wc_sid;                                                        // loopback SID from write command to DID
  ws_hdr[7]  = 1'b1;                                                            // SoT: not supporting fragmentation yet
  ws_hdr[8]  = 1'b1;                                                            // EoT: not supporting fragmentation yet
  ws_hdr[14:9]  = 6'd3;                                                         // Read command
  ws_hdr[17:15]  = wc_did;                                                      // loopback DID from wrtie command to SID
  ws_hdr[19:18]   = wc_id;
end

// declare the state parameters for read
parameter S_RC_HDR = 2'd0;
parameter S_RDS_WAIT = 2'd1;
parameter S_RDS_HDR = 2'd2;
parameter S_RDS_PLD = 2'd3;
assign int_pslverr = 1'd0;
// =======================================================================
// Read Processing
// =======================================================================
// Current Read Flit Count
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rc_cnt <= #1ps 1'd0;
  else if (rc_cnt_en)
    rc_cnt <= #1ps rc_cnt_nxt;
end

assign prdata = int_prdata;
assign pslverr_w = int_pslverr;
// Read State Machine State
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rd_state <= #1ps S_RC_HDR;
  else if (rd_state_en)
    rd_state <= #1ps rd_state_nxt;
end

// Read Command Packing Buffer
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rc_buf[0] <= #1ps {60{1'b0}};
    end
  else
    begin
      if (rc_buf_en[0])
        rc_buf[0] <= #1ps if1_flitdata;
    end
end

assign rc_buf_en = rc_buf_we << rc_cnt;
// ============================================
// Read Data + Status flit sequencer
// ============================================
always_comb
begin
  // Defaults
  rd_state_nxt  = rd_state;
  rc_cnt_nxt    = rc_cnt;
  ir0_req       = 1'b0;
  ir0_sop       = 1'b0;
  ir0_eop       = 1'b0;
  ir0_flitdata  = {34{1'b0}};
  rds_transinfo_we = 1'b0;
  if1_ready     = 1'b0;
  rf_ready      = 1'b0;
  // Write enables
  rd_state_en   = 1'b0;
  rc_cnt_en     = 1'b0;
  rc_buf_we     = 1'b0;
  int_arvalid  = 1'b0;
  case (rd_state)
    S_RC_HDR:
      begin
        if1_ready    = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if1_req)
          begin
            // Header transmission is complete
            if (rc_cnt == 1'd0)
              begin
                int_arvalid  = 1'b1;
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rc_buf_we    = 1'b1;
                rds_transinfo_we = 1'b1;
                rd_state_nxt = S_RDS_WAIT;
                rd_state_en   = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                rc_buf_we    = 1'b1;
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
   S_RDS_WAIT:
   begin
    if (int_pready && int_penable && !int_pwrite)
    begin
        rd_state_nxt = S_RDS_HDR;
        rd_state_en  = 1'b1;
    end
   end
   S_RDS_HDR:
      begin
        ir0_req   = 1'd1;
        ir0_sop   = (rc_cnt == 1'd0);
        case(rc_cnt)
          1'd0: ir0_flitdata = rds_hdr[33:0];
          1'd1: ir0_flitdata = rds_hdr[67:34];
          default: ir0_flitdata = {34{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir0_req && ir0_ready)
          begin
            // Complete header is done
            if (rc_cnt == 1'd1)
              begin
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rd_state_nxt = S_RDS_PLD;
                rd_state_en   = 1'b1;
              end
            else
              begin
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
    S_RDS_PLD:
      begin
        ir0_req       = rf_req;
        ir0_eop       = rf_eop;
        ir0_flitdata  = rf_flitdata;
        rf_ready      = ir0_ready;
        if (rf_req && rf_eop && ir0_ready)
          begin
            rd_state_nxt = S_RC_HDR;
            rd_state_en   = 1'b1;
          end
      end
  endcase
end

always_ff @(posedge rcclk) assert ( (frst_n===1'b0) || (int_arvalid == 1'b0) || (rc_burst != 2'b00) || ({{(32-3){1'b0}},rc_plen} <= (32<<1) ) ) else $error("ERROR usb4_tc_noc_apbtea0 : %0t : Read data burst request is larger than TEA can handle. Read data burst size(rplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,rc_plen,(32<<1) );
usb4_tc_noc_apbtea0_rdpack rdpack (
  .clk(rdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .tr_req(rds_transinfo_we),                                                    // i:1
  .tr_rdy(rds_transinfo_rdy),                                                   // o:1
  .tr_size(rc_size),                                                            // i:3
  .tr_burst(rc_burst),                                                          // i:2
  .tr_addrlsb(rc_addr[11:0]),                                                   // i:12
  .tr_plen(rc_plen),                                                            // i:3
  .r_req(rd_req),                                                               // o:1
  .r_last(rd_last),                                                             // o:1
  .r_data(prdata),                                                              // i:32
  .r_slverr(pslverr_w),                                                         // i:1
  .r_ready(rd_ready),                                                           // i:1
  .f_req(rf_req),                                                               // o:1
  .f_eop(rf_eop),                                                               // o:1
  .f_flitdata(rf_flitdata),                                                     // o:34
  .f_ready(rf_ready),                                                           // i:1
  .tr_addrlsb_out(rc_addr_pack)                                                 // o:12
);
// Create incoming rc bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rc_bus[59:0] = (rd_state == S_RC_HDR) ? if1_flitdata : rc_buf[0];
// assign rc.bus = {$rcBusStr};
// Read Command Signal Unpacking
assign rc_sid = rc_bus[17:15];
assign rc_did = rc_bus[6:4];
assign rc_id = rc_bus[19:18];
assign rc_addr = rc_bus[54:23];
assign rc_qos = rc_bus[3:0];
assign rc_plen = rc_bus[22:20];
assign rc_prot = 3'd0;
assign rc_rawsize = rc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign rc_size = Narrow_Req ? ((rc_rawsize < 3'd2) ? rc_rawsize : 3'd2) : ((rc_rawsize > 3'd2) ? 3'd2 : rc_rawsize);
assign rc_burst = rc_bus[59:58];
assign Narrow_Req = rc_rawsize < 3'd2;
// ============================================
// Read Data + Status Header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  rds_hdr            = {68{1'b0}};
  // Assign over the various fields
  rds_hdr[3:0]  = rc_qos;                                                       // loopback QoS from write command
  rds_hdr[6:4]  = rc_sid;                                                       // loopback SID from write command to DID
  rds_hdr[7]  = 1'b1;                                                           // SoT: not supporting fragmentation yet
  rds_hdr[8]  = 1'b1;                                                           // EoT: not supporting fragmentation yet
  rds_hdr[14:9]  = 6'd1;                                                        // Read data / status
  rds_hdr[17:15]  = rc_did;                                                     // loopback DID from wrtie command to SID
  rds_hdr[19:18]   = rc_id;
  rds_hdr[22:20] = rc_plen;
  rds_hdr[30:23]  = (rc_burst==2'd2) ? 8'(rc_addr[11:0] >> rc_size) : rc_addr[7:0];
  rds_hdr[33:31]  = rc_size;
  rds_hdr[35:34] = rc_burst;
end

// Arbitrate between read and write state machines for use of APB interface
parameter S_PSEL = 2'd0;
parameter S_PWEN = 2'd1;
parameter S_PREN = 2'd2;
parameter S_PRDATA = 2'd3;
// APB State Machine State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_state <= #1ps S_PSEL;
  else if (apb_state_en)
    apb_state <= #1ps apb_state_nxt;
end

// Read / Write Arbiter State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_wrarb <= #1ps 1'd0;
  else if (apb_wrarb_en)
    apb_wrarb <= #1ps apb_wrarb_nxt;
end

// For multiple targets and when both rd and wr are active
always_comb
begin
  int_psel      = 1'b0;
  int_pwrite    = 1'b0;
  int_penable   = 1'b0;
  int_paddr     = {9{1'b0}};
  int_pwdata    = {32{1'b0}};
  int_pstrb     = {4{1'b0}};
  int_pprot     = 3'd0;
  apb_state_nxt = apb_state;
  apb_state_en  = 1'b0;
  apb_wrarb_nxt = apb_wrarb;
  apb_wrarb_en  = 1'b0;
  wr_ready      = 1'b0;
  rd_ready      = 1'b0;
  case (apb_state)
    S_PSEL:
      begin
        if (wr_req && (!rd_req || apb_wrarb))
          begin
            int_psel      = 1'b1;
            int_paddr     = wc_addr_unpack[8:0];
            int_pwrite    = 1'b1;
            int_pwdata    = wr_data;
            int_pstrb     = wr_strb;
            int_pprot     = wc_prot;
            apb_state_nxt = S_PWEN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b0;
            apb_wrarb_en  = 1'b1;
          end
        else if (rd_req)
          begin
            int_psel      = 1'b1;
            int_paddr     = rc_addr_pack[8:0];
            int_pprot     = rc_prot;
            apb_state_nxt = S_PREN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b1;
            apb_wrarb_en  = 1'b1;
          end
      end
    S_PWEN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
        int_pwrite  = 1'b1;
        int_paddr   = wc_addr_unpack[8:0];
        int_pwdata  = wr_data;
        int_pstrb   = wr_strb;
        int_pprot   = wc_prot;
        if (int_pready)
          begin
            wr_ready   = 1'b1;
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
          end
      end
    S_PREN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
            int_paddr     = rc_addr_pack[8:0];
        int_pprot   = rc_prot;
        if (int_pready)
          begin
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
            rd_ready   = 1'b1;
          end
      end
    // S_PRDATA:
    // begin
    // apb.state.nxt = S_PSEL;
    // apb.state.en  = 1'b1;
    // end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_epipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire      [8:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  // dst
  output logic     [8:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata                                             // Read data
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea0_epipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_epipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea0_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea0_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea0_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea0_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_apbcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_wccg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_wdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_f1cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_rdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_wdunpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wtr_req,
  output logic           wtr_rdy,
  input  wire      [2:0] wtr_size,                                              // Transfer size per data phase
  input  wire      [1:0] wtr_burst,                                             // Burst addressing mode
  input  wire     [11:0] wtr_addrlsb,                                           // 12 LSBs of address
  input  wire      [2:0] wtr_plen,                                              // Packet length in bytes
  output logic           w_valid,
  output logic    [31:0] w_data,
  output logic     [3:0] w_strb,
  output logic           w_last,
  input  wire            w_ready,
  input  wire            f_req,
  input  wire            f_eop,
  input  wire     [35:0] f_flitdata,
  output logic           f_ready,
  output logic    [11:0] wtr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [2:0] sizeCnvDiv;
logic     [4:0] firstCnt2Wrap;
logic     [7:0] wtr_mask;
logic     [7:0] wtr_mis;
logic    [10:0] firstXferCnt;
logic    [10:0] xferCnt;
logic    [10:0] xferCnt_nxt;
logic     [0:0] xferCnt_en;
logic    [10:0] useXferCnt;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic    [31:0] muxed_w_data;
logic     [3:0] muxed_w_strb;
logic           flitDone;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic     [0:0] haveFlit;
logic     [0:0] haveFlit_nxt;
logic     [0:0] haveFlit_en;
logic    [35:0] flitData;
logic    [35:0] flitData_nxt;
logic     [0:0] flitData_en;
logic           flitValid;
logic    [11:0] lower_baddr;
logic    [11:0] upper_baddr;
logic    [11:0] lower_addr;
logic    [11:0] upper_addr;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
logic    [11:0] saddr;
logic     [2:0] splen;
// Extracted from packet header
// APB W Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},wtr_plen} - 1'b1;                                    // We only care about 8 bits of address for our word indexing
assign wrapToAddr = wtr_addrlsb[7:0] & ~bamask;                                 // This is the address offset we wrap to
assign wrapIndex = wtr_addrlsb >> wtr_size;
assign sizeCnvDiv = wtr_plen >> wtr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign wtr_mask = (8'b1<<wtr_size) - 1'b1;
assign wtr_mis = wtr_addrlsb[7:0] & wtr_mask;
assign firstXferCnt = (wtr_burst!=2'd1) ? 11'(wtr_plen>>wtr_size) : 11'((16'(wtr_plen)+wtr_mask+wtr_mis)>>wtr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    xferCnt <= #1ps 11'd0;
  else if (xferCnt_en)
    xferCnt <= #1ps xferCnt_nxt;
end

assign useXferCnt = xferCnt;
always_comb
begin
  xferCnt_nxt = xferCnt;
  xferCnt_en  = 1'b0;
  if( newCmd )
    begin
      xferCnt_nxt = firstXferCnt;
      xferCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      xferCnt_nxt = useXferCnt - 1'd1;
      xferCnt_en  = 1'b1;
    end
end

assign wtr_rdy = ~trInPkt;
assign newCmd = wtr_req && wtr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = w_valid && w_ready;
assign f_ready = ~haveFlit || flitDone;
assign w_valid = flitValid;
assign w_last = w_valid && useXferCnt==11'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps wtr_burst;
end

assign use_tr_burst = held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps wtr_size;
end

assign use_tr_size = held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( busWriteValid && w_last )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> wtr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (wtr_addrlsb[7:0] & 8'd3) >> wtr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( w_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone;
assign muxed_w_data[7:0] = flitData[7:0];
assign muxed_w_strb[3:0] = flitData[35:32];
assign muxed_w_data[15:8] = flitData[15:8];
assign muxed_w_data[23:16] = flitData[23:16];
assign muxed_w_data[31:24] = flitData[31:24];
assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    haveFlit <= #1ps 1'd0;
  else if (haveFlit_en)
    haveFlit <= #1ps haveFlit_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitData <= #1ps {36{1'b0}};
  else if (flitData_en)
    flitData <= #1ps flitData_nxt;
end

assign flitValid = haveFlit;
always_comb
begin
  haveFlit_nxt   = haveFlit;
  haveFlit_en    = 1'b0;
  flitData_nxt   = flitData;
  flitData_en    = 1'b0;
  if( flitWriteValid )
    begin
      haveFlit_nxt   = 1'b1;
      haveFlit_en    = 1'b1;
      flitData_en    = 1'b1;
      flitData_nxt   = f_flitdata;
    end
  else if( flitDone )
    begin
      haveFlit_nxt   = 1'b0;
      haveFlit_en    = 1'b1;
    end
end

assign w_data[7:0] = (w_valid && wrMask[0]) ? muxed_w_data[7:0] : 8'd0;
assign w_data[15:8] = (w_valid && wrMask[1]) ? muxed_w_data[15:8] : 8'd0;
assign w_data[23:16] = (w_valid && wrMask[2]) ? muxed_w_data[23:16] : 8'd0;
assign w_data[31:24] = (w_valid && wrMask[3]) ? muxed_w_data[31:24] : 8'd0;
assign w_strb = w_valid ? muxed_w_strb & wrMask : 4'd0;
assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  addrlsb_nxt   = addrlsb;
  // Write enables
  addrlsb_en    = 1'b0;
  if (newCmd)
    begin
      addrlsb_nxt = wtr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred from packing FIFO
  else if (busWriteValid)
    begin
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps wtr_addrlsb;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps wtr_plen;
end

assign wtr_addrlsb_out = !(newCmd) ? addrlsb : wtr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea0_rdpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            tr_req,
  output logic           tr_rdy,
  input  wire      [2:0] tr_size,
  input  wire      [1:0] tr_burst,
  input  wire     [11:0] tr_addrlsb,
  input  wire      [2:0] tr_plen,
  output logic           r_req,
  output logic           r_last,
  input  wire     [31:0] r_data,
  input  wire            r_slverr,
  input  wire            r_ready,
  output logic           f_req,
  output logic           f_eop,
  output logic    [33:0] f_flitdata,
  input  wire            f_ready,
  output logic    [11:0] tr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [4:0] firstCnt2Wrap;
logic     [2:0] sizeCnvDiv;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [0:0] heldFlitDone;
logic     [0:0] heldEop;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isNarrow;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic           flitDone;
logic           useBusWdCnt;
logic    [33:0] flitWd;
logic    [33:0] flitWd_nxt;
logic     [0:0] flitWd_en;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] lower_baddr;                                                    // Lower burst address
logic    [11:0] upper_baddr;                                                    // Upper burst address
logic    [11:0] lower_addr;                                                     // Lower element address
logic    [11:0] upper_addr;                                                     // Upper element address
logic    [11:0] esize_minus_first_offset;
logic    [11:0] first_offset;
logic     [2:0] raw_wcnt;
logic     [2:0] wcnt;
logic    [11:0] saddr;
logic     [2:0] wplen;
logic     [2:0] wplen_nxt;
logic     [0:0] wplen_en;
logic     [2:0] splen;
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
// Extracted from AXI AW Channel
// APB R Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},tr_plen} - 1'b1;                                     // We only care about 8 bits of address for our word indexing
assign wrapToAddr = tr_addrlsb[7:0] & ~bamask;                                  // This is the address offset we wrap to
assign wrapIndex = tr_addrlsb >> tr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign sizeCnvDiv = tr_plen >> tr_size;
assign tr_rdy = ~trInPkt;
assign f_flitdata = flitWd;
assign f_req = heldFlitDone;
assign f_eop = heldEop;
assign r_req = trInPkt_nxt && (!heldFlitDone || flitWriteValid);
assign newCmd = tr_req && tr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = r_ready && r_req;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldFlitDone <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldFlitDone <= #1ps flitDone;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldEop <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldEop <= #1ps flitDone && r_last;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps tr_burst;
end

assign use_tr_burst = (newCmd) ? tr_burst : held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps tr_size;
end

assign use_tr_size = (newCmd) ? tr_size : held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isNarrow = use_tr_size<3'd2;
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( flitWriteValid && f_eop )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> tr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = (newCmd) ? subBusWdCntWrap_nxt : subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = newCmd ? firstCnt2Wrap : cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (tr_addrlsb[7:0] & 8'd3) >> tr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = (newCmd) ? firstSubBusWdCnt[1:0] : subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( r_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone || (isNarrow && busWriteValid);
assign useBusWdCnt = 1'b0;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitWd <= #1ps {34{1'b0}};
  else if (flitWd_en)
    flitWd <= #1ps flitWd_nxt;
end

assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_comb
begin
  // First, assign the bus word to every possible flit word slot
  flitWd_nxt = flitWriteValid ? {34{1'b0}} : flitWd;
  // Start out with nothing enabled
  flitWd_en = flitWriteValid ? 1'b1 : 1'b0;
  // Now enable any bytes that are being written this cycle
  if( busWriteValid )
    begin
      if( useBusWdCnt == 1'd0 )
        begin
          if( wrMask[0] )
            begin
              flitWd_nxt[7:0] = r_data[7:0];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[1] )
            begin
              flitWd_nxt[15:8] = r_data[15:8];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[2] )
            begin
              flitWd_nxt[23:16] = r_data[23:16];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[3] )
            begin
              flitWd_nxt[31:24] = r_data[31:24];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
        end
    end
end

assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
assign esize_minus_first_offset = esize - first_offset;
assign first_offset = addrlsb & amask;
assign raw_wcnt = (held_tr_burst == 2'd1) ? esize_minus_first_offset[2:0] : esize[2:0];
assign wcnt = (raw_wcnt > wplen) ? wplen : raw_wcnt;
assign r_last = (wcnt >= wplen);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps tr_addrlsb;
end

// Write remaining packet length and address LSB tracking flops
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    wplen <= #1ps 3'd0;
  else if (wplen_en)
    wplen <= #1ps wplen_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps tr_plen;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  wplen_nxt   = wplen;
  addrlsb_nxt = addrlsb;
  wplen_en    = 1'b0;
  addrlsb_en  = 1'b0;
  if (tr_req && tr_rdy)
    begin
      wplen_nxt   = tr_plen;
      wplen_en    = 1'b1;
      addrlsb_nxt = tr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred to packing FIFO
  else if (busWriteValid)
    begin
      wplen_en    = 1'b1;
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            wplen_nxt   = wplen - wcnt;
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            wplen_nxt   = wplen   - wcnt;
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            wplen_nxt   = wplen      - wcnt;
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            wplen_nxt   = wplen;
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

assign tr_addrlsb_out = !(newCmd) ? addrlsb : tr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1 (
  input  wire            clk,
  input  wire            rst_n,
  // t
  output logic    [15:0] t_paddr,                                               // Address
  output logic           t_psel,                                                // Select
  output logic           t_penable,                                             // Enable
  output logic           t_pwrite,                                              // Write not read
  output logic    [31:0] t_pwdata,                                              // Write data
  output logic     [3:0] t_pstrb,                                               // Write strobes
  input  wire            t_pready,                                              // Ready
  input  wire     [31:0] t_prdata,                                              // Read data
  // f0
  input  wire            f0_activity,                                           // Upcoming activity indicator
  input  wire            f0_req,                                                // Flit transfer request
  input  wire            f0_sop,                                                // Start of packet indicator
  input  wire            f0_eop,                                                // End of packet indicator
  input  wire     [35:0] f0_flitdata,                                           // Flit data
  output logic           f0_ready,                                              // Flit transfer ready
  // f1
  input  wire            f1_activity,                                           // Upcoming activity indicator
  input  wire            f1_req,                                                // Flit transfer request
  input  wire            f1_sop,                                                // Start of packet indicator
  input  wire            f1_eop,                                                // End of packet indicator
  input  wire     [59:0] f1_flitdata,                                           // Flit data
  output logic           f1_ready,                                              // Flit transfer ready
  // r0
  output logic           r0_activity,                                           // Upcoming activity indicator
  output logic           r0_req,                                                // Flit transfer request
  output logic           r0_sop,                                                // Start of packet indicator
  output logic           r0_eop,                                                // End of packet indicator
  output logic    [33:0] r0_flitdata,                                           // Flit data
  input  wire            r0_ready,                                              // Flit transfer ready
  // r1
  output logic           r1_activity,                                           // Upcoming activity indicator
  output logic           r1_req,                                                // Flit transfer request
  output logic           r1_sop,                                                // Start of packet indicator
  output logic           r1_eop,                                                // End of packet indicator
  output logic    [23:0] r1_flitdata,                                           // Flit data
  input  wire            r1_ready                                               // Flit transfer ready
);

logic    [15:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic           wr_req;
logic           wr_ready;
logic           wr_last;
logic    [31:0] wr_data;
logic     [3:0] wr_strb;
logic           wc_buf_we;
logic    [71:0] wc_bus;
logic     [2:0] wc_sid;
logic     [2:0] wc_did;
logic     [1:0] wc_id;
logic    [31:0] wc_addr;
logic     [7:0] wc_len;
logic     [2:0] wc_rawsize;
logic     [2:0] wc_size;
logic     [1:0] wc_burst;
logic     [3:0] wc_qos;
logic     [2:0] wc_plen;
logic     [2:0] wc_prot;
logic           wcd_transinfo_en;
logic           wcd_transinfo_rdy;
logic           wf_req;
logic           wf_eop;
logic    [35:0] wf_flitdata;
logic           wf_ready;
logic    [23:0] ws_hdr;
logic           int_awvalid;
logic    [67:0] rds_hdr;
logic           rd_req;
logic           rd_ready;
logic           rd_last;
logic           rc_buf_we;
logic    [59:0] rc_bus;
logic     [2:0] rc_sid;
logic     [2:0] rc_did;
logic     [1:0] rc_id;
logic    [31:0] rc_addr;
logic     [2:0] rc_rawsize;
logic     [2:0] rc_size;
logic     [1:0] rc_burst;
logic     [3:0] rc_qos;
logic     [2:0] rc_plen;
logic     [2:0] rc_prot;
logic           rf_req;
logic           rf_eop;
logic    [33:0] rf_flitdata;
logic           rf_ready;
logic           rds_transinfo_we;
logic           rds_transinfo_rdy;
logic           int_arvalid;
logic    [11:0] wc_addr_unpack;
logic    [11:0] rc_addr_pack;
logic     [2:0] int_pprot;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           apbclk;
logic           apbclkAct;
logic           int_apbactivity;
logic           wcclk;
logic           wcclkAct;
wire            int_awactivity;
logic           wdclk;
logic           wdclkAct;
logic           int_wactivity;
logic           rcclk;
logic           rcclkAct;
logic           int_aractivity;
logic           rdclk;
logic           rdclkAct;
logic           rdclkEn;
logic           wrDone;
logic     [0:0] wr_cnt;
logic     [0:0] wr_cnt_nxt;
logic     [0:0] wr_cnt_en;
logic     [1:0] wr_state;
logic     [1:0] wr_state_nxt;
logic     [0:0] wr_state_en;
logic    [35:0] wc_buf [1:0];
logic     [1:0] wc_buf_en;
logic           int_pslverr;
logic     [0:0] rc_cnt;
logic     [0:0] rc_cnt_nxt;
logic     [0:0] rc_cnt_en;
logic           pslverr_w;
logic    [31:0] prdata;
logic     [1:0] rd_state;
logic     [1:0] rd_state_nxt;
logic     [0:0] rd_state_en;
logic    [59:0] rc_buf [0:0];
logic     [0:0] rc_buf_en;
logic           Narrow_Req;
logic     [1:0] apb_state;
logic     [1:0] apb_state_nxt;
logic     [0:0] apb_state_en;
logic     [0:0] apb_wrarb;
logic     [0:0] apb_wrarb_nxt;
logic     [0:0] apb_wrarb_en;
// ========================================================================//
// Parameter Declarations
// ========================================================================//
// ========================================================================//
// Process parameters and create local derived variables
// ========================================================================//
// ========================================================================//
// Define module I/O
// ========================================================================//
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Target Interface(s) (APB manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Egress APB Pipeline Component
usb4_tc_noc_apbtea1_epipe epipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(int_paddr),                                                        // i:16
  .src_psel(int_psel),                                                          // i:1
  .src_penable(int_penable),                                                    // i:1
  .src_pwrite(int_pwrite),                                                      // i:1
  .src_pwdata(int_pwdata),                                                      // i:32
  .src_pstrb(int_pstrb),                                                        // i:4
  .src_pready(int_pready),                                                      // o:1
  .src_prdata(int_prdata),                                                      // o:32
  .dst_paddr(t_paddr),                                                          // o:16
  .dst_psel(t_psel),                                                            // o:1
  .dst_penable(t_penable),                                                      // o:1
  .dst_pwrite(t_pwrite),                                                        // o:1
  .dst_pwdata(t_pwdata),                                                        // o:32
  .dst_pstrb(t_pstrb),                                                          // o:4
  .dst_pready(t_pready),                                                        // i:1
  .dst_prdata(t_prdata)                                                         // i:32
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea1_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f0_activity),                                                   // i:1
  .src_req(f0_req),                                                             // i:1
  .src_sop(f0_sop),                                                             // i:1
  .src_eop(f0_eop),                                                             // i:1
  .src_flitdata(f0_flitdata),                                                   // i:36
  .src_ready(f0_ready),                                                         // o:1
  .dst_activity(if0_activity),                                                  // o:1
  .dst_req(if0_req),                                                            // o:1
  .dst_sop(if0_sop),                                                            // o:1
  .dst_eop(if0_eop),                                                            // o:1
  .dst_flitdata(if0_flitdata),                                                  // o:36
  .dst_ready(if0_ready)                                                         // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea1_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f1_activity),                                                   // i:1
  .src_req(f1_req),                                                             // i:1
  .src_sop(f1_sop),                                                             // i:1
  .src_eop(f1_eop),                                                             // i:1
  .src_flitdata(f1_flitdata),                                                   // i:60
  .src_ready(f1_ready),                                                         // o:1
  .dst_activity(if1_activity),                                                  // o:1
  .dst_req(if1_req),                                                            // o:1
  .dst_sop(if1_sop),                                                            // o:1
  .dst_eop(if1_eop),                                                            // o:1
  .dst_flitdata(if1_flitdata),                                                  // o:60
  .dst_ready(if1_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea1_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir0_activity),                                                  // i:1
  .src_req(ir0_req),                                                            // i:1
  .src_sop(ir0_sop),                                                            // i:1
  .src_eop(ir0_eop),                                                            // i:1
  .src_flitdata(ir0_flitdata),                                                  // i:34
  .src_ready(ir0_ready),                                                        // o:1
  .dst_activity(r0_activity),                                                   // o:1
  .dst_req(r0_req),                                                             // o:1
  .dst_sop(r0_sop),                                                             // o:1
  .dst_eop(r0_eop),                                                             // o:1
  .dst_flitdata(r0_flitdata),                                                   // o:34
  .dst_ready(r0_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea1_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir1_activity),                                                  // i:1
  .src_req(ir1_req),                                                            // i:1
  .src_sop(ir1_sop),                                                            // i:1
  .src_eop(ir1_eop),                                                            // i:1
  .src_flitdata(ir1_flitdata),                                                  // i:24
  .src_ready(ir1_ready),                                                        // o:1
  .dst_activity(r1_activity),                                                   // o:1
  .dst_req(r1_req),                                                             // o:1
  .dst_sop(r1_sop),                                                             // o:1
  .dst_eop(r1_eop),                                                             // o:1
  .dst_flitdata(r1_flitdata),                                                   // o:24
  .dst_ready(r1_ready)                                                          // i:1
);
// =======================================================================
// Signal declarations
// =======================================================================
// Write Command + Data Sequencer Signals
// Write Command Signals
// Write Response Fields
// Read Data + Status fields
// Read Data + Status Flit Sequencer Signals
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea1_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign int_apbactivity = int_awactivity || int_aractivity;
usb4_tc_noc_apbtea1_apbcg apbcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_apbactivity),                                                      // i:1
  .clkOut(apbclk),                                                              // o:1
  .isActive(apbclkAct)                                                          // o:1
);
assign int_awactivity = if0_activity || if0_req || int_awvalid || ir1_req || wr_req;
usb4_tc_noc_apbtea1_wccg wccg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_awactivity),                                                       // i:1
  .clkOut(wcclk),                                                               // o:1
  .isActive(wcclkAct)                                                           // o:1
);
assign int_wactivity = if0_activity || if0_req || !wcd_transinfo_rdy || int_awvalid;
usb4_tc_noc_apbtea1_wdcg wdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_wactivity),                                                        // i:1
  .clkOut(wdclk),                                                               // o:1
  .isActive(wdclkAct)                                                           // o:1
);
assign ir1_activity = ir1_req;
assign int_aractivity = if1_activity || if1_req || ir0_req || rd_req;
usb4_tc_noc_apbtea1_f1cg f1cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_aractivity),                                                       // i:1
  .clkOut(rcclk),                                                               // o:1
  .isActive(rcclkAct)                                                           // o:1
);
assign ir0_activity = ir0_req;
assign rdclkEn = ir0_activity || if1_activity || if1_req || !rds_transinfo_rdy;
usb4_tc_noc_apbtea1_rdcg rdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(rdclkEn),                                                              // i:1
  .clkOut(rdclk),                                                               // o:1
  .isActive(rdclkAct)                                                           // o:1
);
// =======================================================================
// Write Processing
// =======================================================================
assign wrDone = wr_last && int_penable && int_pwrite && int_pready;
parameter S_WR_HDR = 2'd0;
parameter S_WR_DATA = 2'd1;
parameter S_WR_WAIT = 2'd2;
parameter S_WR_STS = 2'd3;
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign wc_bus[35:0] = wc_buf[0];
assign wc_bus[71:36] = ((wr_state == 2'b00) && (wr_cnt >= 1'd1)) ? if0_flitdata : wc_buf[1];
// Current Flit Count
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_cnt <= #1ps 1'd0;
  else if (wr_cnt_en)
    wr_cnt <= #1ps wr_cnt_nxt;
end

// Write State Machine State
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_state <= #1ps S_WR_HDR;
  else if (wr_state_en)
    wr_state <= #1ps wr_state_nxt;
end

// Write Command Packing Buffer
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      wc_buf[0] <= #1ps {36{1'b0}};
      wc_buf[1] <= #1ps {36{1'b0}};
    end
  else
    begin
      if (wc_buf_en[0])
        wc_buf[0] <= #1ps if0_flitdata;
      if (wc_buf_en[1])
        wc_buf[1] <= #1ps if0_flitdata;
    end
end

assign wc_buf_en = wc_buf_we << wr_cnt;
always_comb
begin
  // Defaults
  if0_ready    = 1'b0;
  ir1_req      = 1'b0;
  ir1_sop      = 1'b0;
  ir1_eop      = 1'b0;
  ir1_flitdata = {24{1'b0}};
  wr_cnt_nxt   = wr_cnt;
  wr_state_nxt = wr_state;
  wcd_transinfo_en = 1'b0;
  wf_req       = 1'b0;
  wf_eop       = 1'b0;
  wf_flitdata  = {36{1'b0}};
  // Write enables
  wc_buf_we    = 1'b0;
  wr_cnt_en    = 1'b0;
  wr_state_en  = 1'b0;
  int_awvalid   = 1'b0;
  case (wr_state)
    S_WR_HDR:
      begin
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_req)
          begin
            if0_ready    = 1'b1;
            // Header transmission is complete
            if (wr_cnt == 1'd1)
              begin
                int_awvalid = wcd_transinfo_rdy;
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wc_buf_we    = 1'b1;
                wcd_transinfo_en = 1'b1;
                wr_state_nxt = S_WR_DATA;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
                wc_buf_we  = 1'b1;
              end
          end
      end
   S_WR_DATA:
      begin
        wf_req      = if0_req;
        wf_eop      = if0_eop;
        wf_flitdata = if0_flitdata;
        if0_ready   = wf_ready;
        if (if0_req && wf_ready && if0_eop)
          begin
            wr_state_nxt = S_WR_WAIT;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_WAIT:
      begin
        if (wr_req && wr_ready && wr_last)
          begin
            wr_state_nxt = S_WR_STS;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_STS:
      begin
        ir1_req   = 1'b1;
        ir1_sop   = (wr_cnt == 1'd0);
        ir1_eop   = (wr_cnt == 1'd0);
        case(wr_cnt)
          1'd0: ir1_flitdata = ws_hdr[23:0];
          default: ir1_flitdata = {24{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_ready)
          begin
            // Header transmission is complete
            if (wr_cnt == 1'd0)
              begin
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wr_state_nxt = S_WR_HDR;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
              end
          end
      end
  endcase
end

 always_ff @(posedge wcclk) assert ( (frst_n===1'b0) || (int_awvalid == 1'b0) || (wc_burst != 2'b00) || ( {{(32-3){1'b0}},wc_plen} <= (32<<1) )) else $error("ERROR usb4_tc_noc_apbtea1 : %0t : Write data burst request is larger than TEA can handle. Write data burst size(wplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,wc_plen,(32<<1) );
usb4_tc_noc_apbtea1_wdunpack wdunpack (
  .clk(wdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .wtr_req(wcd_transinfo_en),                                                   // i:1
  .wtr_rdy(wcd_transinfo_rdy),                                                  // o:1
  .wtr_size(wc_size),                                                           // i:3
  .wtr_burst(wc_burst),                                                         // i:2
  .wtr_addrlsb(wc_addr[11:0]),                                                  // i:12
  .wtr_plen(wc_plen),                                                           // i:3
  .w_valid(wr_req),                                                             // o:1
  .w_data(wr_data),                                                             // o:32
  .w_strb(wr_strb),                                                             // o:4
  .w_last(wr_last),                                                             // o:1
  .w_ready(wr_ready),                                                           // i:1
  .f_req(wf_req),                                                               // i:1
  .f_eop(wf_eop),                                                               // i:1
  .f_flitdata(wf_flitdata),                                                     // i:36
  .f_ready(wf_ready),                                                           // o:1
  .wtr_addrlsb_out(wc_addr_unpack)                                              // o:12
);
// Write Command + Data Signal Unpacking
assign wc_sid = wc_bus[17:15];
assign wc_did = wc_bus[6:4];
assign wc_id = wc_bus[19:18];
assign wc_addr = wc_bus[54:23];
assign wc_qos = wc_bus[3:0];
assign wc_plen = wc_bus[22:20];
assign wc_prot = 3'd0;
assign wc_rawsize = wc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign wc_size = (wc_rawsize > 3'd2) ? 3'd2 : wc_rawsize;
assign wc_burst = wc_bus[59:58];
// =======================================================================
// Write Response Path Processing
// =======================================================================
// ============================================
// Write Response header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  ws_hdr            = {24{1'b0}};
  // Assign over the various fields
  ws_hdr[3:0]  = wc_qos;                                                        // loopback QoS from write command
  ws_hdr[6:4]  = wc_sid;                                                        // loopback SID from write command to DID
  ws_hdr[7]  = 1'b1;                                                            // SoT: not supporting fragmentation yet
  ws_hdr[8]  = 1'b1;                                                            // EoT: not supporting fragmentation yet
  ws_hdr[14:9]  = 6'd3;                                                         // Read command
  ws_hdr[17:15]  = wc_did;                                                      // loopback DID from wrtie command to SID
  ws_hdr[19:18]   = wc_id;
end

// declare the state parameters for read
parameter S_RC_HDR = 2'd0;
parameter S_RDS_WAIT = 2'd1;
parameter S_RDS_HDR = 2'd2;
parameter S_RDS_PLD = 2'd3;
assign int_pslverr = 1'd0;
// =======================================================================
// Read Processing
// =======================================================================
// Current Read Flit Count
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rc_cnt <= #1ps 1'd0;
  else if (rc_cnt_en)
    rc_cnt <= #1ps rc_cnt_nxt;
end

assign prdata = int_prdata;
assign pslverr_w = int_pslverr;
// Read State Machine State
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rd_state <= #1ps S_RC_HDR;
  else if (rd_state_en)
    rd_state <= #1ps rd_state_nxt;
end

// Read Command Packing Buffer
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rc_buf[0] <= #1ps {60{1'b0}};
    end
  else
    begin
      if (rc_buf_en[0])
        rc_buf[0] <= #1ps if1_flitdata;
    end
end

assign rc_buf_en = rc_buf_we << rc_cnt;
// ============================================
// Read Data + Status flit sequencer
// ============================================
always_comb
begin
  // Defaults
  rd_state_nxt  = rd_state;
  rc_cnt_nxt    = rc_cnt;
  ir0_req       = 1'b0;
  ir0_sop       = 1'b0;
  ir0_eop       = 1'b0;
  ir0_flitdata  = {34{1'b0}};
  rds_transinfo_we = 1'b0;
  if1_ready     = 1'b0;
  rf_ready      = 1'b0;
  // Write enables
  rd_state_en   = 1'b0;
  rc_cnt_en     = 1'b0;
  rc_buf_we     = 1'b0;
  int_arvalid  = 1'b0;
  case (rd_state)
    S_RC_HDR:
      begin
        if1_ready    = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if1_req)
          begin
            // Header transmission is complete
            if (rc_cnt == 1'd0)
              begin
                int_arvalid  = 1'b1;
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rc_buf_we    = 1'b1;
                rds_transinfo_we = 1'b1;
                rd_state_nxt = S_RDS_WAIT;
                rd_state_en   = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                rc_buf_we    = 1'b1;
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
   S_RDS_WAIT:
   begin
    if (int_pready && int_penable && !int_pwrite)
    begin
        rd_state_nxt = S_RDS_HDR;
        rd_state_en  = 1'b1;
    end
   end
   S_RDS_HDR:
      begin
        ir0_req   = 1'd1;
        ir0_sop   = (rc_cnt == 1'd0);
        case(rc_cnt)
          1'd0: ir0_flitdata = rds_hdr[33:0];
          1'd1: ir0_flitdata = rds_hdr[67:34];
          default: ir0_flitdata = {34{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir0_req && ir0_ready)
          begin
            // Complete header is done
            if (rc_cnt == 1'd1)
              begin
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rd_state_nxt = S_RDS_PLD;
                rd_state_en   = 1'b1;
              end
            else
              begin
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
    S_RDS_PLD:
      begin
        ir0_req       = rf_req;
        ir0_eop       = rf_eop;
        ir0_flitdata  = rf_flitdata;
        rf_ready      = ir0_ready;
        if (rf_req && rf_eop && ir0_ready)
          begin
            rd_state_nxt = S_RC_HDR;
            rd_state_en   = 1'b1;
          end
      end
  endcase
end

always_ff @(posedge rcclk) assert ( (frst_n===1'b0) || (int_arvalid == 1'b0) || (rc_burst != 2'b00) || ({{(32-3){1'b0}},rc_plen} <= (32<<1) ) ) else $error("ERROR usb4_tc_noc_apbtea1 : %0t : Read data burst request is larger than TEA can handle. Read data burst size(rplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,rc_plen,(32<<1) );
usb4_tc_noc_apbtea1_rdpack rdpack (
  .clk(rdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .tr_req(rds_transinfo_we),                                                    // i:1
  .tr_rdy(rds_transinfo_rdy),                                                   // o:1
  .tr_size(rc_size),                                                            // i:3
  .tr_burst(rc_burst),                                                          // i:2
  .tr_addrlsb(rc_addr[11:0]),                                                   // i:12
  .tr_plen(rc_plen),                                                            // i:3
  .r_req(rd_req),                                                               // o:1
  .r_last(rd_last),                                                             // o:1
  .r_data(prdata),                                                              // i:32
  .r_slverr(pslverr_w),                                                         // i:1
  .r_ready(rd_ready),                                                           // i:1
  .f_req(rf_req),                                                               // o:1
  .f_eop(rf_eop),                                                               // o:1
  .f_flitdata(rf_flitdata),                                                     // o:34
  .f_ready(rf_ready),                                                           // i:1
  .tr_addrlsb_out(rc_addr_pack)                                                 // o:12
);
// Create incoming rc bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rc_bus[59:0] = (rd_state == S_RC_HDR) ? if1_flitdata : rc_buf[0];
// assign rc.bus = {$rcBusStr};
// Read Command Signal Unpacking
assign rc_sid = rc_bus[17:15];
assign rc_did = rc_bus[6:4];
assign rc_id = rc_bus[19:18];
assign rc_addr = rc_bus[54:23];
assign rc_qos = rc_bus[3:0];
assign rc_plen = rc_bus[22:20];
assign rc_prot = 3'd0;
assign rc_rawsize = rc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign rc_size = Narrow_Req ? ((rc_rawsize < 3'd2) ? rc_rawsize : 3'd2) : ((rc_rawsize > 3'd2) ? 3'd2 : rc_rawsize);
assign rc_burst = rc_bus[59:58];
assign Narrow_Req = rc_rawsize < 3'd2;
// ============================================
// Read Data + Status Header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  rds_hdr            = {68{1'b0}};
  // Assign over the various fields
  rds_hdr[3:0]  = rc_qos;                                                       // loopback QoS from write command
  rds_hdr[6:4]  = rc_sid;                                                       // loopback SID from write command to DID
  rds_hdr[7]  = 1'b1;                                                           // SoT: not supporting fragmentation yet
  rds_hdr[8]  = 1'b1;                                                           // EoT: not supporting fragmentation yet
  rds_hdr[14:9]  = 6'd1;                                                        // Read data / status
  rds_hdr[17:15]  = rc_did;                                                     // loopback DID from wrtie command to SID
  rds_hdr[19:18]   = rc_id;
  rds_hdr[22:20] = rc_plen;
  rds_hdr[30:23]  = (rc_burst==2'd2) ? 8'(rc_addr[11:0] >> rc_size) : rc_addr[7:0];
  rds_hdr[33:31]  = rc_size;
  rds_hdr[35:34] = rc_burst;
end

// Arbitrate between read and write state machines for use of APB interface
parameter S_PSEL = 2'd0;
parameter S_PWEN = 2'd1;
parameter S_PREN = 2'd2;
parameter S_PRDATA = 2'd3;
// APB State Machine State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_state <= #1ps S_PSEL;
  else if (apb_state_en)
    apb_state <= #1ps apb_state_nxt;
end

// Read / Write Arbiter State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_wrarb <= #1ps 1'd0;
  else if (apb_wrarb_en)
    apb_wrarb <= #1ps apb_wrarb_nxt;
end

// For multiple targets and when both rd and wr are active
always_comb
begin
  int_psel      = 1'b0;
  int_pwrite    = 1'b0;
  int_penable   = 1'b0;
  int_paddr     = {16{1'b0}};
  int_pwdata    = {32{1'b0}};
  int_pstrb     = {4{1'b0}};
  int_pprot     = 3'd0;
  apb_state_nxt = apb_state;
  apb_state_en  = 1'b0;
  apb_wrarb_nxt = apb_wrarb;
  apb_wrarb_en  = 1'b0;
  wr_ready      = 1'b0;
  rd_ready      = 1'b0;
  case (apb_state)
    S_PSEL:
      begin
        if (wr_req && (!rd_req || apb_wrarb))
          begin
            int_psel      = 1'b1;
            int_paddr     = {wc_addr[15:12],wc_addr_unpack};
            int_pwrite    = 1'b1;
            int_pwdata    = wr_data;
            int_pstrb     = wr_strb;
            int_pprot     = wc_prot;
            apb_state_nxt = S_PWEN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b0;
            apb_wrarb_en  = 1'b1;
          end
        else if (rd_req)
          begin
            int_psel      = 1'b1;
            int_paddr     = {rc_addr[15:12],rc_addr_pack};
            int_pprot     = rc_prot;
            apb_state_nxt = S_PREN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b1;
            apb_wrarb_en  = 1'b1;
          end
      end
    S_PWEN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
        int_pwrite  = 1'b1;
        int_paddr   = {wc_addr[15:12],wc_addr_unpack};
        int_pwdata  = wr_data;
        int_pstrb   = wr_strb;
        int_pprot   = wc_prot;
        if (int_pready)
          begin
            wr_ready   = 1'b1;
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
          end
      end
    S_PREN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
            int_paddr     = {rc_addr[15:12],rc_addr_pack};
        int_pprot   = rc_prot;
        if (int_pready)
          begin
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
            rd_ready   = 1'b1;
          end
      end
    // S_PRDATA:
    // begin
    // apb.state.nxt = S_PSEL;
    // apb.state.en  = 1'b1;
    // end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_epipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire     [15:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  // dst
  output logic    [15:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata                                             // Read data
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea1_epipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_epipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea1_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea1_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea1_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea1_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_apbcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_wccg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_wdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_f1cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_rdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_wdunpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wtr_req,
  output logic           wtr_rdy,
  input  wire      [2:0] wtr_size,                                              // Transfer size per data phase
  input  wire      [1:0] wtr_burst,                                             // Burst addressing mode
  input  wire     [11:0] wtr_addrlsb,                                           // 12 LSBs of address
  input  wire      [2:0] wtr_plen,                                              // Packet length in bytes
  output logic           w_valid,
  output logic    [31:0] w_data,
  output logic     [3:0] w_strb,
  output logic           w_last,
  input  wire            w_ready,
  input  wire            f_req,
  input  wire            f_eop,
  input  wire     [35:0] f_flitdata,
  output logic           f_ready,
  output logic    [11:0] wtr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [2:0] sizeCnvDiv;
logic     [4:0] firstCnt2Wrap;
logic     [7:0] wtr_mask;
logic     [7:0] wtr_mis;
logic    [10:0] firstXferCnt;
logic    [10:0] xferCnt;
logic    [10:0] xferCnt_nxt;
logic     [0:0] xferCnt_en;
logic    [10:0] useXferCnt;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic    [31:0] muxed_w_data;
logic     [3:0] muxed_w_strb;
logic           flitDone;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic     [0:0] haveFlit;
logic     [0:0] haveFlit_nxt;
logic     [0:0] haveFlit_en;
logic    [35:0] flitData;
logic    [35:0] flitData_nxt;
logic     [0:0] flitData_en;
logic           flitValid;
logic    [11:0] lower_baddr;
logic    [11:0] upper_baddr;
logic    [11:0] lower_addr;
logic    [11:0] upper_addr;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
logic    [11:0] saddr;
logic     [2:0] splen;
// Extracted from packet header
// APB W Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},wtr_plen} - 1'b1;                                    // We only care about 8 bits of address for our word indexing
assign wrapToAddr = wtr_addrlsb[7:0] & ~bamask;                                 // This is the address offset we wrap to
assign wrapIndex = wtr_addrlsb >> wtr_size;
assign sizeCnvDiv = wtr_plen >> wtr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign wtr_mask = (8'b1<<wtr_size) - 1'b1;
assign wtr_mis = wtr_addrlsb[7:0] & wtr_mask;
assign firstXferCnt = (wtr_burst!=2'd1) ? 11'(wtr_plen>>wtr_size) : 11'((16'(wtr_plen)+wtr_mask+wtr_mis)>>wtr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    xferCnt <= #1ps 11'd0;
  else if (xferCnt_en)
    xferCnt <= #1ps xferCnt_nxt;
end

assign useXferCnt = xferCnt;
always_comb
begin
  xferCnt_nxt = xferCnt;
  xferCnt_en  = 1'b0;
  if( newCmd )
    begin
      xferCnt_nxt = firstXferCnt;
      xferCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      xferCnt_nxt = useXferCnt - 1'd1;
      xferCnt_en  = 1'b1;
    end
end

assign wtr_rdy = ~trInPkt;
assign newCmd = wtr_req && wtr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = w_valid && w_ready;
assign f_ready = ~haveFlit || flitDone;
assign w_valid = flitValid;
assign w_last = w_valid && useXferCnt==11'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps wtr_burst;
end

assign use_tr_burst = held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps wtr_size;
end

assign use_tr_size = held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( busWriteValid && w_last )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> wtr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (wtr_addrlsb[7:0] & 8'd3) >> wtr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( w_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone;
assign muxed_w_data[7:0] = flitData[7:0];
assign muxed_w_strb[3:0] = flitData[35:32];
assign muxed_w_data[15:8] = flitData[15:8];
assign muxed_w_data[23:16] = flitData[23:16];
assign muxed_w_data[31:24] = flitData[31:24];
assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    haveFlit <= #1ps 1'd0;
  else if (haveFlit_en)
    haveFlit <= #1ps haveFlit_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitData <= #1ps {36{1'b0}};
  else if (flitData_en)
    flitData <= #1ps flitData_nxt;
end

assign flitValid = haveFlit;
always_comb
begin
  haveFlit_nxt   = haveFlit;
  haveFlit_en    = 1'b0;
  flitData_nxt   = flitData;
  flitData_en    = 1'b0;
  if( flitWriteValid )
    begin
      haveFlit_nxt   = 1'b1;
      haveFlit_en    = 1'b1;
      flitData_en    = 1'b1;
      flitData_nxt   = f_flitdata;
    end
  else if( flitDone )
    begin
      haveFlit_nxt   = 1'b0;
      haveFlit_en    = 1'b1;
    end
end

assign w_data[7:0] = (w_valid && wrMask[0]) ? muxed_w_data[7:0] : 8'd0;
assign w_data[15:8] = (w_valid && wrMask[1]) ? muxed_w_data[15:8] : 8'd0;
assign w_data[23:16] = (w_valid && wrMask[2]) ? muxed_w_data[23:16] : 8'd0;
assign w_data[31:24] = (w_valid && wrMask[3]) ? muxed_w_data[31:24] : 8'd0;
assign w_strb = w_valid ? muxed_w_strb & wrMask : 4'd0;
assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  addrlsb_nxt   = addrlsb;
  // Write enables
  addrlsb_en    = 1'b0;
  if (newCmd)
    begin
      addrlsb_nxt = wtr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred from packing FIFO
  else if (busWriteValid)
    begin
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps wtr_addrlsb;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps wtr_plen;
end

assign wtr_addrlsb_out = !(newCmd) ? addrlsb : wtr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea1_rdpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            tr_req,
  output logic           tr_rdy,
  input  wire      [2:0] tr_size,
  input  wire      [1:0] tr_burst,
  input  wire     [11:0] tr_addrlsb,
  input  wire      [2:0] tr_plen,
  output logic           r_req,
  output logic           r_last,
  input  wire     [31:0] r_data,
  input  wire            r_slverr,
  input  wire            r_ready,
  output logic           f_req,
  output logic           f_eop,
  output logic    [33:0] f_flitdata,
  input  wire            f_ready,
  output logic    [11:0] tr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [4:0] firstCnt2Wrap;
logic     [2:0] sizeCnvDiv;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [0:0] heldFlitDone;
logic     [0:0] heldEop;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isNarrow;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic           flitDone;
logic           useBusWdCnt;
logic    [33:0] flitWd;
logic    [33:0] flitWd_nxt;
logic     [0:0] flitWd_en;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] lower_baddr;                                                    // Lower burst address
logic    [11:0] upper_baddr;                                                    // Upper burst address
logic    [11:0] lower_addr;                                                     // Lower element address
logic    [11:0] upper_addr;                                                     // Upper element address
logic    [11:0] esize_minus_first_offset;
logic    [11:0] first_offset;
logic     [2:0] raw_wcnt;
logic     [2:0] wcnt;
logic    [11:0] saddr;
logic     [2:0] wplen;
logic     [2:0] wplen_nxt;
logic     [0:0] wplen_en;
logic     [2:0] splen;
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
// Extracted from AXI AW Channel
// APB R Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},tr_plen} - 1'b1;                                     // We only care about 8 bits of address for our word indexing
assign wrapToAddr = tr_addrlsb[7:0] & ~bamask;                                  // This is the address offset we wrap to
assign wrapIndex = tr_addrlsb >> tr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign sizeCnvDiv = tr_plen >> tr_size;
assign tr_rdy = ~trInPkt;
assign f_flitdata = flitWd;
assign f_req = heldFlitDone;
assign f_eop = heldEop;
assign r_req = trInPkt_nxt && (!heldFlitDone || flitWriteValid);
assign newCmd = tr_req && tr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = r_ready && r_req;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldFlitDone <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldFlitDone <= #1ps flitDone;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldEop <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldEop <= #1ps flitDone && r_last;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps tr_burst;
end

assign use_tr_burst = (newCmd) ? tr_burst : held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps tr_size;
end

assign use_tr_size = (newCmd) ? tr_size : held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isNarrow = use_tr_size<3'd2;
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( flitWriteValid && f_eop )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> tr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = (newCmd) ? subBusWdCntWrap_nxt : subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = newCmd ? firstCnt2Wrap : cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (tr_addrlsb[7:0] & 8'd3) >> tr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = (newCmd) ? firstSubBusWdCnt[1:0] : subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( r_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone || (isNarrow && busWriteValid);
assign useBusWdCnt = 1'b0;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitWd <= #1ps {34{1'b0}};
  else if (flitWd_en)
    flitWd <= #1ps flitWd_nxt;
end

assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_comb
begin
  // First, assign the bus word to every possible flit word slot
  flitWd_nxt = flitWriteValid ? {34{1'b0}} : flitWd;
  // Start out with nothing enabled
  flitWd_en = flitWriteValid ? 1'b1 : 1'b0;
  // Now enable any bytes that are being written this cycle
  if( busWriteValid )
    begin
      if( useBusWdCnt == 1'd0 )
        begin
          if( wrMask[0] )
            begin
              flitWd_nxt[7:0] = r_data[7:0];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[1] )
            begin
              flitWd_nxt[15:8] = r_data[15:8];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[2] )
            begin
              flitWd_nxt[23:16] = r_data[23:16];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[3] )
            begin
              flitWd_nxt[31:24] = r_data[31:24];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
        end
    end
end

assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
assign esize_minus_first_offset = esize - first_offset;
assign first_offset = addrlsb & amask;
assign raw_wcnt = (held_tr_burst == 2'd1) ? esize_minus_first_offset[2:0] : esize[2:0];
assign wcnt = (raw_wcnt > wplen) ? wplen : raw_wcnt;
assign r_last = (wcnt >= wplen);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps tr_addrlsb;
end

// Write remaining packet length and address LSB tracking flops
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    wplen <= #1ps 3'd0;
  else if (wplen_en)
    wplen <= #1ps wplen_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps tr_plen;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  wplen_nxt   = wplen;
  addrlsb_nxt = addrlsb;
  wplen_en    = 1'b0;
  addrlsb_en  = 1'b0;
  if (tr_req && tr_rdy)
    begin
      wplen_nxt   = tr_plen;
      wplen_en    = 1'b1;
      addrlsb_nxt = tr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred to packing FIFO
  else if (busWriteValid)
    begin
      wplen_en    = 1'b1;
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            wplen_nxt   = wplen - wcnt;
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            wplen_nxt   = wplen   - wcnt;
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            wplen_nxt   = wplen      - wcnt;
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            wplen_nxt   = wplen;
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

assign tr_addrlsb_out = !(newCmd) ? addrlsb : tr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2 (
  input  wire            clk,
  input  wire            rst_n,
  // t
  output logic    [15:0] t_paddr,                                               // Address
  output logic           t_psel,                                                // Select
  output logic           t_penable,                                             // Enable
  output logic           t_pwrite,                                              // Write not read
  output logic    [31:0] t_pwdata,                                              // Write data
  output logic     [3:0] t_pstrb,                                               // Write strobes
  input  wire            t_pready,                                              // Ready
  input  wire     [31:0] t_prdata,                                              // Read data
  // f0
  input  wire            f0_activity,                                           // Upcoming activity indicator
  input  wire            f0_req,                                                // Flit transfer request
  input  wire            f0_sop,                                                // Start of packet indicator
  input  wire            f0_eop,                                                // End of packet indicator
  input  wire     [35:0] f0_flitdata,                                           // Flit data
  output logic           f0_ready,                                              // Flit transfer ready
  // f1
  input  wire            f1_activity,                                           // Upcoming activity indicator
  input  wire            f1_req,                                                // Flit transfer request
  input  wire            f1_sop,                                                // Start of packet indicator
  input  wire            f1_eop,                                                // End of packet indicator
  input  wire     [59:0] f1_flitdata,                                           // Flit data
  output logic           f1_ready,                                              // Flit transfer ready
  // r0
  output logic           r0_activity,                                           // Upcoming activity indicator
  output logic           r0_req,                                                // Flit transfer request
  output logic           r0_sop,                                                // Start of packet indicator
  output logic           r0_eop,                                                // End of packet indicator
  output logic    [33:0] r0_flitdata,                                           // Flit data
  input  wire            r0_ready,                                              // Flit transfer ready
  // r1
  output logic           r1_activity,                                           // Upcoming activity indicator
  output logic           r1_req,                                                // Flit transfer request
  output logic           r1_sop,                                                // Start of packet indicator
  output logic           r1_eop,                                                // End of packet indicator
  output logic    [23:0] r1_flitdata,                                           // Flit data
  input  wire            r1_ready                                               // Flit transfer ready
);

logic    [15:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic           wr_req;
logic           wr_ready;
logic           wr_last;
logic    [31:0] wr_data;
logic     [3:0] wr_strb;
logic           wc_buf_we;
logic    [71:0] wc_bus;
logic     [2:0] wc_sid;
logic     [2:0] wc_did;
logic     [1:0] wc_id;
logic    [31:0] wc_addr;
logic     [7:0] wc_len;
logic     [2:0] wc_rawsize;
logic     [2:0] wc_size;
logic     [1:0] wc_burst;
logic     [3:0] wc_qos;
logic     [2:0] wc_plen;
logic     [2:0] wc_prot;
logic           wcd_transinfo_en;
logic           wcd_transinfo_rdy;
logic           wf_req;
logic           wf_eop;
logic    [35:0] wf_flitdata;
logic           wf_ready;
logic    [23:0] ws_hdr;
logic           int_awvalid;
logic    [67:0] rds_hdr;
logic           rd_req;
logic           rd_ready;
logic           rd_last;
logic           rc_buf_we;
logic    [59:0] rc_bus;
logic     [2:0] rc_sid;
logic     [2:0] rc_did;
logic     [1:0] rc_id;
logic    [31:0] rc_addr;
logic     [2:0] rc_rawsize;
logic     [2:0] rc_size;
logic     [1:0] rc_burst;
logic     [3:0] rc_qos;
logic     [2:0] rc_plen;
logic     [2:0] rc_prot;
logic           rf_req;
logic           rf_eop;
logic    [33:0] rf_flitdata;
logic           rf_ready;
logic           rds_transinfo_we;
logic           rds_transinfo_rdy;
logic           int_arvalid;
logic    [11:0] wc_addr_unpack;
logic    [11:0] rc_addr_pack;
logic     [2:0] int_pprot;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           apbclk;
logic           apbclkAct;
logic           int_apbactivity;
logic           wcclk;
logic           wcclkAct;
wire            int_awactivity;
logic           wdclk;
logic           wdclkAct;
logic           int_wactivity;
logic           rcclk;
logic           rcclkAct;
logic           int_aractivity;
logic           rdclk;
logic           rdclkAct;
logic           rdclkEn;
logic           wrDone;
logic     [0:0] wr_cnt;
logic     [0:0] wr_cnt_nxt;
logic     [0:0] wr_cnt_en;
logic     [1:0] wr_state;
logic     [1:0] wr_state_nxt;
logic     [0:0] wr_state_en;
logic    [35:0] wc_buf [1:0];
logic     [1:0] wc_buf_en;
logic           int_pslverr;
logic     [0:0] rc_cnt;
logic     [0:0] rc_cnt_nxt;
logic     [0:0] rc_cnt_en;
logic           pslverr_w;
logic    [31:0] prdata;
logic     [1:0] rd_state;
logic     [1:0] rd_state_nxt;
logic     [0:0] rd_state_en;
logic    [59:0] rc_buf [0:0];
logic     [0:0] rc_buf_en;
logic           Narrow_Req;
logic     [1:0] apb_state;
logic     [1:0] apb_state_nxt;
logic     [0:0] apb_state_en;
logic     [0:0] apb_wrarb;
logic     [0:0] apb_wrarb_nxt;
logic     [0:0] apb_wrarb_en;
// ========================================================================//
// Parameter Declarations
// ========================================================================//
// ========================================================================//
// Process parameters and create local derived variables
// ========================================================================//
// ========================================================================//
// Define module I/O
// ========================================================================//
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Target Interface(s) (APB manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Egress APB Pipeline Component
usb4_tc_noc_apbtea2_epipe epipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(int_paddr),                                                        // i:16
  .src_psel(int_psel),                                                          // i:1
  .src_penable(int_penable),                                                    // i:1
  .src_pwrite(int_pwrite),                                                      // i:1
  .src_pwdata(int_pwdata),                                                      // i:32
  .src_pstrb(int_pstrb),                                                        // i:4
  .src_pready(int_pready),                                                      // o:1
  .src_prdata(int_prdata),                                                      // o:32
  .dst_paddr(t_paddr),                                                          // o:16
  .dst_psel(t_psel),                                                            // o:1
  .dst_penable(t_penable),                                                      // o:1
  .dst_pwrite(t_pwrite),                                                        // o:1
  .dst_pwdata(t_pwdata),                                                        // o:32
  .dst_pstrb(t_pstrb),                                                          // o:4
  .dst_pready(t_pready),                                                        // i:1
  .dst_prdata(t_prdata)                                                         // i:32
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea2_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f0_activity),                                                   // i:1
  .src_req(f0_req),                                                             // i:1
  .src_sop(f0_sop),                                                             // i:1
  .src_eop(f0_eop),                                                             // i:1
  .src_flitdata(f0_flitdata),                                                   // i:36
  .src_ready(f0_ready),                                                         // o:1
  .dst_activity(if0_activity),                                                  // o:1
  .dst_req(if0_req),                                                            // o:1
  .dst_sop(if0_sop),                                                            // o:1
  .dst_eop(if0_eop),                                                            // o:1
  .dst_flitdata(if0_flitdata),                                                  // o:36
  .dst_ready(if0_ready)                                                         // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea2_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f1_activity),                                                   // i:1
  .src_req(f1_req),                                                             // i:1
  .src_sop(f1_sop),                                                             // i:1
  .src_eop(f1_eop),                                                             // i:1
  .src_flitdata(f1_flitdata),                                                   // i:60
  .src_ready(f1_ready),                                                         // o:1
  .dst_activity(if1_activity),                                                  // o:1
  .dst_req(if1_req),                                                            // o:1
  .dst_sop(if1_sop),                                                            // o:1
  .dst_eop(if1_eop),                                                            // o:1
  .dst_flitdata(if1_flitdata),                                                  // o:60
  .dst_ready(if1_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea2_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir0_activity),                                                  // i:1
  .src_req(ir0_req),                                                            // i:1
  .src_sop(ir0_sop),                                                            // i:1
  .src_eop(ir0_eop),                                                            // i:1
  .src_flitdata(ir0_flitdata),                                                  // i:34
  .src_ready(ir0_ready),                                                        // o:1
  .dst_activity(r0_activity),                                                   // o:1
  .dst_req(r0_req),                                                             // o:1
  .dst_sop(r0_sop),                                                             // o:1
  .dst_eop(r0_eop),                                                             // o:1
  .dst_flitdata(r0_flitdata),                                                   // o:34
  .dst_ready(r0_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea2_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir1_activity),                                                  // i:1
  .src_req(ir1_req),                                                            // i:1
  .src_sop(ir1_sop),                                                            // i:1
  .src_eop(ir1_eop),                                                            // i:1
  .src_flitdata(ir1_flitdata),                                                  // i:24
  .src_ready(ir1_ready),                                                        // o:1
  .dst_activity(r1_activity),                                                   // o:1
  .dst_req(r1_req),                                                             // o:1
  .dst_sop(r1_sop),                                                             // o:1
  .dst_eop(r1_eop),                                                             // o:1
  .dst_flitdata(r1_flitdata),                                                   // o:24
  .dst_ready(r1_ready)                                                          // i:1
);
// =======================================================================
// Signal declarations
// =======================================================================
// Write Command + Data Sequencer Signals
// Write Command Signals
// Write Response Fields
// Read Data + Status fields
// Read Data + Status Flit Sequencer Signals
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea2_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign int_apbactivity = int_awactivity || int_aractivity;
usb4_tc_noc_apbtea2_apbcg apbcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_apbactivity),                                                      // i:1
  .clkOut(apbclk),                                                              // o:1
  .isActive(apbclkAct)                                                          // o:1
);
assign int_awactivity = if0_activity || if0_req || int_awvalid || ir1_req || wr_req;
usb4_tc_noc_apbtea2_wccg wccg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_awactivity),                                                       // i:1
  .clkOut(wcclk),                                                               // o:1
  .isActive(wcclkAct)                                                           // o:1
);
assign int_wactivity = if0_activity || if0_req || !wcd_transinfo_rdy || int_awvalid;
usb4_tc_noc_apbtea2_wdcg wdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_wactivity),                                                        // i:1
  .clkOut(wdclk),                                                               // o:1
  .isActive(wdclkAct)                                                           // o:1
);
assign ir1_activity = ir1_req;
assign int_aractivity = if1_activity || if1_req || ir0_req || rd_req;
usb4_tc_noc_apbtea2_f1cg f1cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_aractivity),                                                       // i:1
  .clkOut(rcclk),                                                               // o:1
  .isActive(rcclkAct)                                                           // o:1
);
assign ir0_activity = ir0_req;
assign rdclkEn = ir0_activity || if1_activity || if1_req || !rds_transinfo_rdy;
usb4_tc_noc_apbtea2_rdcg rdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(rdclkEn),                                                              // i:1
  .clkOut(rdclk),                                                               // o:1
  .isActive(rdclkAct)                                                           // o:1
);
// =======================================================================
// Write Processing
// =======================================================================
assign wrDone = wr_last && int_penable && int_pwrite && int_pready;
parameter S_WR_HDR = 2'd0;
parameter S_WR_DATA = 2'd1;
parameter S_WR_WAIT = 2'd2;
parameter S_WR_STS = 2'd3;
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign wc_bus[35:0] = wc_buf[0];
assign wc_bus[71:36] = ((wr_state == 2'b00) && (wr_cnt >= 1'd1)) ? if0_flitdata : wc_buf[1];
// Current Flit Count
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_cnt <= #1ps 1'd0;
  else if (wr_cnt_en)
    wr_cnt <= #1ps wr_cnt_nxt;
end

// Write State Machine State
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_state <= #1ps S_WR_HDR;
  else if (wr_state_en)
    wr_state <= #1ps wr_state_nxt;
end

// Write Command Packing Buffer
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      wc_buf[0] <= #1ps {36{1'b0}};
      wc_buf[1] <= #1ps {36{1'b0}};
    end
  else
    begin
      if (wc_buf_en[0])
        wc_buf[0] <= #1ps if0_flitdata;
      if (wc_buf_en[1])
        wc_buf[1] <= #1ps if0_flitdata;
    end
end

assign wc_buf_en = wc_buf_we << wr_cnt;
always_comb
begin
  // Defaults
  if0_ready    = 1'b0;
  ir1_req      = 1'b0;
  ir1_sop      = 1'b0;
  ir1_eop      = 1'b0;
  ir1_flitdata = {24{1'b0}};
  wr_cnt_nxt   = wr_cnt;
  wr_state_nxt = wr_state;
  wcd_transinfo_en = 1'b0;
  wf_req       = 1'b0;
  wf_eop       = 1'b0;
  wf_flitdata  = {36{1'b0}};
  // Write enables
  wc_buf_we    = 1'b0;
  wr_cnt_en    = 1'b0;
  wr_state_en  = 1'b0;
  int_awvalid   = 1'b0;
  case (wr_state)
    S_WR_HDR:
      begin
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_req)
          begin
            if0_ready    = 1'b1;
            // Header transmission is complete
            if (wr_cnt == 1'd1)
              begin
                int_awvalid = wcd_transinfo_rdy;
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wc_buf_we    = 1'b1;
                wcd_transinfo_en = 1'b1;
                wr_state_nxt = S_WR_DATA;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
                wc_buf_we  = 1'b1;
              end
          end
      end
   S_WR_DATA:
      begin
        wf_req      = if0_req;
        wf_eop      = if0_eop;
        wf_flitdata = if0_flitdata;
        if0_ready   = wf_ready;
        if (if0_req && wf_ready && if0_eop)
          begin
            wr_state_nxt = S_WR_WAIT;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_WAIT:
      begin
        if (wr_req && wr_ready && wr_last)
          begin
            wr_state_nxt = S_WR_STS;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_STS:
      begin
        ir1_req   = 1'b1;
        ir1_sop   = (wr_cnt == 1'd0);
        ir1_eop   = (wr_cnt == 1'd0);
        case(wr_cnt)
          1'd0: ir1_flitdata = ws_hdr[23:0];
          default: ir1_flitdata = {24{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_ready)
          begin
            // Header transmission is complete
            if (wr_cnt == 1'd0)
              begin
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wr_state_nxt = S_WR_HDR;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
              end
          end
      end
  endcase
end

 always_ff @(posedge wcclk) assert ( (frst_n===1'b0) || (int_awvalid == 1'b0) || (wc_burst != 2'b00) || ( {{(32-3){1'b0}},wc_plen} <= (32<<1) )) else $error("ERROR usb4_tc_noc_apbtea2 : %0t : Write data burst request is larger than TEA can handle. Write data burst size(wplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,wc_plen,(32<<1) );
usb4_tc_noc_apbtea2_wdunpack wdunpack (
  .clk(wdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .wtr_req(wcd_transinfo_en),                                                   // i:1
  .wtr_rdy(wcd_transinfo_rdy),                                                  // o:1
  .wtr_size(wc_size),                                                           // i:3
  .wtr_burst(wc_burst),                                                         // i:2
  .wtr_addrlsb(wc_addr[11:0]),                                                  // i:12
  .wtr_plen(wc_plen),                                                           // i:3
  .w_valid(wr_req),                                                             // o:1
  .w_data(wr_data),                                                             // o:32
  .w_strb(wr_strb),                                                             // o:4
  .w_last(wr_last),                                                             // o:1
  .w_ready(wr_ready),                                                           // i:1
  .f_req(wf_req),                                                               // i:1
  .f_eop(wf_eop),                                                               // i:1
  .f_flitdata(wf_flitdata),                                                     // i:36
  .f_ready(wf_ready),                                                           // o:1
  .wtr_addrlsb_out(wc_addr_unpack)                                              // o:12
);
// Write Command + Data Signal Unpacking
assign wc_sid = wc_bus[17:15];
assign wc_did = wc_bus[6:4];
assign wc_id = wc_bus[19:18];
assign wc_addr = wc_bus[54:23];
assign wc_qos = wc_bus[3:0];
assign wc_plen = wc_bus[22:20];
assign wc_prot = 3'd0;
assign wc_rawsize = wc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign wc_size = (wc_rawsize > 3'd2) ? 3'd2 : wc_rawsize;
assign wc_burst = wc_bus[59:58];
// =======================================================================
// Write Response Path Processing
// =======================================================================
// ============================================
// Write Response header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  ws_hdr            = {24{1'b0}};
  // Assign over the various fields
  ws_hdr[3:0]  = wc_qos;                                                        // loopback QoS from write command
  ws_hdr[6:4]  = wc_sid;                                                        // loopback SID from write command to DID
  ws_hdr[7]  = 1'b1;                                                            // SoT: not supporting fragmentation yet
  ws_hdr[8]  = 1'b1;                                                            // EoT: not supporting fragmentation yet
  ws_hdr[14:9]  = 6'd3;                                                         // Read command
  ws_hdr[17:15]  = wc_did;                                                      // loopback DID from wrtie command to SID
  ws_hdr[19:18]   = wc_id;
end

// declare the state parameters for read
parameter S_RC_HDR = 2'd0;
parameter S_RDS_WAIT = 2'd1;
parameter S_RDS_HDR = 2'd2;
parameter S_RDS_PLD = 2'd3;
assign int_pslverr = 1'd0;
// =======================================================================
// Read Processing
// =======================================================================
// Current Read Flit Count
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rc_cnt <= #1ps 1'd0;
  else if (rc_cnt_en)
    rc_cnt <= #1ps rc_cnt_nxt;
end

assign prdata = int_prdata;
assign pslverr_w = int_pslverr;
// Read State Machine State
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rd_state <= #1ps S_RC_HDR;
  else if (rd_state_en)
    rd_state <= #1ps rd_state_nxt;
end

// Read Command Packing Buffer
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rc_buf[0] <= #1ps {60{1'b0}};
    end
  else
    begin
      if (rc_buf_en[0])
        rc_buf[0] <= #1ps if1_flitdata;
    end
end

assign rc_buf_en = rc_buf_we << rc_cnt;
// ============================================
// Read Data + Status flit sequencer
// ============================================
always_comb
begin
  // Defaults
  rd_state_nxt  = rd_state;
  rc_cnt_nxt    = rc_cnt;
  ir0_req       = 1'b0;
  ir0_sop       = 1'b0;
  ir0_eop       = 1'b0;
  ir0_flitdata  = {34{1'b0}};
  rds_transinfo_we = 1'b0;
  if1_ready     = 1'b0;
  rf_ready      = 1'b0;
  // Write enables
  rd_state_en   = 1'b0;
  rc_cnt_en     = 1'b0;
  rc_buf_we     = 1'b0;
  int_arvalid  = 1'b0;
  case (rd_state)
    S_RC_HDR:
      begin
        if1_ready    = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if1_req)
          begin
            // Header transmission is complete
            if (rc_cnt == 1'd0)
              begin
                int_arvalid  = 1'b1;
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rc_buf_we    = 1'b1;
                rds_transinfo_we = 1'b1;
                rd_state_nxt = S_RDS_WAIT;
                rd_state_en   = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                rc_buf_we    = 1'b1;
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
   S_RDS_WAIT:
   begin
    if (int_pready && int_penable && !int_pwrite)
    begin
        rd_state_nxt = S_RDS_HDR;
        rd_state_en  = 1'b1;
    end
   end
   S_RDS_HDR:
      begin
        ir0_req   = 1'd1;
        ir0_sop   = (rc_cnt == 1'd0);
        case(rc_cnt)
          1'd0: ir0_flitdata = rds_hdr[33:0];
          1'd1: ir0_flitdata = rds_hdr[67:34];
          default: ir0_flitdata = {34{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir0_req && ir0_ready)
          begin
            // Complete header is done
            if (rc_cnt == 1'd1)
              begin
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rd_state_nxt = S_RDS_PLD;
                rd_state_en   = 1'b1;
              end
            else
              begin
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
    S_RDS_PLD:
      begin
        ir0_req       = rf_req;
        ir0_eop       = rf_eop;
        ir0_flitdata  = rf_flitdata;
        rf_ready      = ir0_ready;
        if (rf_req && rf_eop && ir0_ready)
          begin
            rd_state_nxt = S_RC_HDR;
            rd_state_en   = 1'b1;
          end
      end
  endcase
end

always_ff @(posedge rcclk) assert ( (frst_n===1'b0) || (int_arvalid == 1'b0) || (rc_burst != 2'b00) || ({{(32-3){1'b0}},rc_plen} <= (32<<1) ) ) else $error("ERROR usb4_tc_noc_apbtea2 : %0t : Read data burst request is larger than TEA can handle. Read data burst size(rplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,rc_plen,(32<<1) );
usb4_tc_noc_apbtea2_rdpack rdpack (
  .clk(rdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .tr_req(rds_transinfo_we),                                                    // i:1
  .tr_rdy(rds_transinfo_rdy),                                                   // o:1
  .tr_size(rc_size),                                                            // i:3
  .tr_burst(rc_burst),                                                          // i:2
  .tr_addrlsb(rc_addr[11:0]),                                                   // i:12
  .tr_plen(rc_plen),                                                            // i:3
  .r_req(rd_req),                                                               // o:1
  .r_last(rd_last),                                                             // o:1
  .r_data(prdata),                                                              // i:32
  .r_slverr(pslverr_w),                                                         // i:1
  .r_ready(rd_ready),                                                           // i:1
  .f_req(rf_req),                                                               // o:1
  .f_eop(rf_eop),                                                               // o:1
  .f_flitdata(rf_flitdata),                                                     // o:34
  .f_ready(rf_ready),                                                           // i:1
  .tr_addrlsb_out(rc_addr_pack)                                                 // o:12
);
// Create incoming rc bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rc_bus[59:0] = (rd_state == S_RC_HDR) ? if1_flitdata : rc_buf[0];
// assign rc.bus = {$rcBusStr};
// Read Command Signal Unpacking
assign rc_sid = rc_bus[17:15];
assign rc_did = rc_bus[6:4];
assign rc_id = rc_bus[19:18];
assign rc_addr = rc_bus[54:23];
assign rc_qos = rc_bus[3:0];
assign rc_plen = rc_bus[22:20];
assign rc_prot = 3'd0;
assign rc_rawsize = rc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign rc_size = Narrow_Req ? ((rc_rawsize < 3'd2) ? rc_rawsize : 3'd2) : ((rc_rawsize > 3'd2) ? 3'd2 : rc_rawsize);
assign rc_burst = rc_bus[59:58];
assign Narrow_Req = rc_rawsize < 3'd2;
// ============================================
// Read Data + Status Header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  rds_hdr            = {68{1'b0}};
  // Assign over the various fields
  rds_hdr[3:0]  = rc_qos;                                                       // loopback QoS from write command
  rds_hdr[6:4]  = rc_sid;                                                       // loopback SID from write command to DID
  rds_hdr[7]  = 1'b1;                                                           // SoT: not supporting fragmentation yet
  rds_hdr[8]  = 1'b1;                                                           // EoT: not supporting fragmentation yet
  rds_hdr[14:9]  = 6'd1;                                                        // Read data / status
  rds_hdr[17:15]  = rc_did;                                                     // loopback DID from wrtie command to SID
  rds_hdr[19:18]   = rc_id;
  rds_hdr[22:20] = rc_plen;
  rds_hdr[30:23]  = (rc_burst==2'd2) ? 8'(rc_addr[11:0] >> rc_size) : rc_addr[7:0];
  rds_hdr[33:31]  = rc_size;
  rds_hdr[35:34] = rc_burst;
end

// Arbitrate between read and write state machines for use of APB interface
parameter S_PSEL = 2'd0;
parameter S_PWEN = 2'd1;
parameter S_PREN = 2'd2;
parameter S_PRDATA = 2'd3;
// APB State Machine State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_state <= #1ps S_PSEL;
  else if (apb_state_en)
    apb_state <= #1ps apb_state_nxt;
end

// Read / Write Arbiter State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_wrarb <= #1ps 1'd0;
  else if (apb_wrarb_en)
    apb_wrarb <= #1ps apb_wrarb_nxt;
end

// For multiple targets and when both rd and wr are active
always_comb
begin
  int_psel      = 1'b0;
  int_pwrite    = 1'b0;
  int_penable   = 1'b0;
  int_paddr     = {16{1'b0}};
  int_pwdata    = {32{1'b0}};
  int_pstrb     = {4{1'b0}};
  int_pprot     = 3'd0;
  apb_state_nxt = apb_state;
  apb_state_en  = 1'b0;
  apb_wrarb_nxt = apb_wrarb;
  apb_wrarb_en  = 1'b0;
  wr_ready      = 1'b0;
  rd_ready      = 1'b0;
  case (apb_state)
    S_PSEL:
      begin
        if (wr_req && (!rd_req || apb_wrarb))
          begin
            int_psel      = 1'b1;
            int_paddr     = {wc_addr[15:12],wc_addr_unpack};
            int_pwrite    = 1'b1;
            int_pwdata    = wr_data;
            int_pstrb     = wr_strb;
            int_pprot     = wc_prot;
            apb_state_nxt = S_PWEN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b0;
            apb_wrarb_en  = 1'b1;
          end
        else if (rd_req)
          begin
            int_psel      = 1'b1;
            int_paddr     = {rc_addr[15:12],rc_addr_pack};
            int_pprot     = rc_prot;
            apb_state_nxt = S_PREN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b1;
            apb_wrarb_en  = 1'b1;
          end
      end
    S_PWEN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
        int_pwrite  = 1'b1;
        int_paddr   = {wc_addr[15:12],wc_addr_unpack};
        int_pwdata  = wr_data;
        int_pstrb   = wr_strb;
        int_pprot   = wc_prot;
        if (int_pready)
          begin
            wr_ready   = 1'b1;
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
          end
      end
    S_PREN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
            int_paddr     = {rc_addr[15:12],rc_addr_pack};
        int_pprot   = rc_prot;
        if (int_pready)
          begin
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
            rd_ready   = 1'b1;
          end
      end
    // S_PRDATA:
    // begin
    // apb.state.nxt = S_PSEL;
    // apb.state.en  = 1'b1;
    // end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_epipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire     [15:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  // dst
  output logic    [15:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata                                             // Read data
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea2_epipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_epipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea2_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea2_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea2_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea2_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_apbcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_wccg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_wdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_f1cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_rdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_wdunpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wtr_req,
  output logic           wtr_rdy,
  input  wire      [2:0] wtr_size,                                              // Transfer size per data phase
  input  wire      [1:0] wtr_burst,                                             // Burst addressing mode
  input  wire     [11:0] wtr_addrlsb,                                           // 12 LSBs of address
  input  wire      [2:0] wtr_plen,                                              // Packet length in bytes
  output logic           w_valid,
  output logic    [31:0] w_data,
  output logic     [3:0] w_strb,
  output logic           w_last,
  input  wire            w_ready,
  input  wire            f_req,
  input  wire            f_eop,
  input  wire     [35:0] f_flitdata,
  output logic           f_ready,
  output logic    [11:0] wtr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [2:0] sizeCnvDiv;
logic     [4:0] firstCnt2Wrap;
logic     [7:0] wtr_mask;
logic     [7:0] wtr_mis;
logic    [10:0] firstXferCnt;
logic    [10:0] xferCnt;
logic    [10:0] xferCnt_nxt;
logic     [0:0] xferCnt_en;
logic    [10:0] useXferCnt;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic    [31:0] muxed_w_data;
logic     [3:0] muxed_w_strb;
logic           flitDone;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic     [0:0] haveFlit;
logic     [0:0] haveFlit_nxt;
logic     [0:0] haveFlit_en;
logic    [35:0] flitData;
logic    [35:0] flitData_nxt;
logic     [0:0] flitData_en;
logic           flitValid;
logic    [11:0] lower_baddr;
logic    [11:0] upper_baddr;
logic    [11:0] lower_addr;
logic    [11:0] upper_addr;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
logic    [11:0] saddr;
logic     [2:0] splen;
// Extracted from packet header
// APB W Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},wtr_plen} - 1'b1;                                    // We only care about 8 bits of address for our word indexing
assign wrapToAddr = wtr_addrlsb[7:0] & ~bamask;                                 // This is the address offset we wrap to
assign wrapIndex = wtr_addrlsb >> wtr_size;
assign sizeCnvDiv = wtr_plen >> wtr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign wtr_mask = (8'b1<<wtr_size) - 1'b1;
assign wtr_mis = wtr_addrlsb[7:0] & wtr_mask;
assign firstXferCnt = (wtr_burst!=2'd1) ? 11'(wtr_plen>>wtr_size) : 11'((16'(wtr_plen)+wtr_mask+wtr_mis)>>wtr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    xferCnt <= #1ps 11'd0;
  else if (xferCnt_en)
    xferCnt <= #1ps xferCnt_nxt;
end

assign useXferCnt = xferCnt;
always_comb
begin
  xferCnt_nxt = xferCnt;
  xferCnt_en  = 1'b0;
  if( newCmd )
    begin
      xferCnt_nxt = firstXferCnt;
      xferCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      xferCnt_nxt = useXferCnt - 1'd1;
      xferCnt_en  = 1'b1;
    end
end

assign wtr_rdy = ~trInPkt;
assign newCmd = wtr_req && wtr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = w_valid && w_ready;
assign f_ready = ~haveFlit || flitDone;
assign w_valid = flitValid;
assign w_last = w_valid && useXferCnt==11'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps wtr_burst;
end

assign use_tr_burst = held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps wtr_size;
end

assign use_tr_size = held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( busWriteValid && w_last )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> wtr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (wtr_addrlsb[7:0] & 8'd3) >> wtr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( w_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone;
assign muxed_w_data[7:0] = flitData[7:0];
assign muxed_w_strb[3:0] = flitData[35:32];
assign muxed_w_data[15:8] = flitData[15:8];
assign muxed_w_data[23:16] = flitData[23:16];
assign muxed_w_data[31:24] = flitData[31:24];
assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    haveFlit <= #1ps 1'd0;
  else if (haveFlit_en)
    haveFlit <= #1ps haveFlit_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitData <= #1ps {36{1'b0}};
  else if (flitData_en)
    flitData <= #1ps flitData_nxt;
end

assign flitValid = haveFlit;
always_comb
begin
  haveFlit_nxt   = haveFlit;
  haveFlit_en    = 1'b0;
  flitData_nxt   = flitData;
  flitData_en    = 1'b0;
  if( flitWriteValid )
    begin
      haveFlit_nxt   = 1'b1;
      haveFlit_en    = 1'b1;
      flitData_en    = 1'b1;
      flitData_nxt   = f_flitdata;
    end
  else if( flitDone )
    begin
      haveFlit_nxt   = 1'b0;
      haveFlit_en    = 1'b1;
    end
end

assign w_data[7:0] = (w_valid && wrMask[0]) ? muxed_w_data[7:0] : 8'd0;
assign w_data[15:8] = (w_valid && wrMask[1]) ? muxed_w_data[15:8] : 8'd0;
assign w_data[23:16] = (w_valid && wrMask[2]) ? muxed_w_data[23:16] : 8'd0;
assign w_data[31:24] = (w_valid && wrMask[3]) ? muxed_w_data[31:24] : 8'd0;
assign w_strb = w_valid ? muxed_w_strb & wrMask : 4'd0;
assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  addrlsb_nxt   = addrlsb;
  // Write enables
  addrlsb_en    = 1'b0;
  if (newCmd)
    begin
      addrlsb_nxt = wtr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred from packing FIFO
  else if (busWriteValid)
    begin
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps wtr_addrlsb;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps wtr_plen;
end

assign wtr_addrlsb_out = !(newCmd) ? addrlsb : wtr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea2_rdpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            tr_req,
  output logic           tr_rdy,
  input  wire      [2:0] tr_size,
  input  wire      [1:0] tr_burst,
  input  wire     [11:0] tr_addrlsb,
  input  wire      [2:0] tr_plen,
  output logic           r_req,
  output logic           r_last,
  input  wire     [31:0] r_data,
  input  wire            r_slverr,
  input  wire            r_ready,
  output logic           f_req,
  output logic           f_eop,
  output logic    [33:0] f_flitdata,
  input  wire            f_ready,
  output logic    [11:0] tr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [4:0] firstCnt2Wrap;
logic     [2:0] sizeCnvDiv;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [0:0] heldFlitDone;
logic     [0:0] heldEop;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isNarrow;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic           flitDone;
logic           useBusWdCnt;
logic    [33:0] flitWd;
logic    [33:0] flitWd_nxt;
logic     [0:0] flitWd_en;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] lower_baddr;                                                    // Lower burst address
logic    [11:0] upper_baddr;                                                    // Upper burst address
logic    [11:0] lower_addr;                                                     // Lower element address
logic    [11:0] upper_addr;                                                     // Upper element address
logic    [11:0] esize_minus_first_offset;
logic    [11:0] first_offset;
logic     [2:0] raw_wcnt;
logic     [2:0] wcnt;
logic    [11:0] saddr;
logic     [2:0] wplen;
logic     [2:0] wplen_nxt;
logic     [0:0] wplen_en;
logic     [2:0] splen;
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
// Extracted from AXI AW Channel
// APB R Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},tr_plen} - 1'b1;                                     // We only care about 8 bits of address for our word indexing
assign wrapToAddr = tr_addrlsb[7:0] & ~bamask;                                  // This is the address offset we wrap to
assign wrapIndex = tr_addrlsb >> tr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign sizeCnvDiv = tr_plen >> tr_size;
assign tr_rdy = ~trInPkt;
assign f_flitdata = flitWd;
assign f_req = heldFlitDone;
assign f_eop = heldEop;
assign r_req = trInPkt_nxt && (!heldFlitDone || flitWriteValid);
assign newCmd = tr_req && tr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = r_ready && r_req;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldFlitDone <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldFlitDone <= #1ps flitDone;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldEop <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldEop <= #1ps flitDone && r_last;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps tr_burst;
end

assign use_tr_burst = (newCmd) ? tr_burst : held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps tr_size;
end

assign use_tr_size = (newCmd) ? tr_size : held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isNarrow = use_tr_size<3'd2;
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( flitWriteValid && f_eop )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> tr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = (newCmd) ? subBusWdCntWrap_nxt : subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = newCmd ? firstCnt2Wrap : cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (tr_addrlsb[7:0] & 8'd3) >> tr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = (newCmd) ? firstSubBusWdCnt[1:0] : subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( r_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone || (isNarrow && busWriteValid);
assign useBusWdCnt = 1'b0;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitWd <= #1ps {34{1'b0}};
  else if (flitWd_en)
    flitWd <= #1ps flitWd_nxt;
end

assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_comb
begin
  // First, assign the bus word to every possible flit word slot
  flitWd_nxt = flitWriteValid ? {34{1'b0}} : flitWd;
  // Start out with nothing enabled
  flitWd_en = flitWriteValid ? 1'b1 : 1'b0;
  // Now enable any bytes that are being written this cycle
  if( busWriteValid )
    begin
      if( useBusWdCnt == 1'd0 )
        begin
          if( wrMask[0] )
            begin
              flitWd_nxt[7:0] = r_data[7:0];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[1] )
            begin
              flitWd_nxt[15:8] = r_data[15:8];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[2] )
            begin
              flitWd_nxt[23:16] = r_data[23:16];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[3] )
            begin
              flitWd_nxt[31:24] = r_data[31:24];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
        end
    end
end

assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
assign esize_minus_first_offset = esize - first_offset;
assign first_offset = addrlsb & amask;
assign raw_wcnt = (held_tr_burst == 2'd1) ? esize_minus_first_offset[2:0] : esize[2:0];
assign wcnt = (raw_wcnt > wplen) ? wplen : raw_wcnt;
assign r_last = (wcnt >= wplen);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps tr_addrlsb;
end

// Write remaining packet length and address LSB tracking flops
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    wplen <= #1ps 3'd0;
  else if (wplen_en)
    wplen <= #1ps wplen_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps tr_plen;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  wplen_nxt   = wplen;
  addrlsb_nxt = addrlsb;
  wplen_en    = 1'b0;
  addrlsb_en  = 1'b0;
  if (tr_req && tr_rdy)
    begin
      wplen_nxt   = tr_plen;
      wplen_en    = 1'b1;
      addrlsb_nxt = tr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred to packing FIFO
  else if (busWriteValid)
    begin
      wplen_en    = 1'b1;
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            wplen_nxt   = wplen - wcnt;
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            wplen_nxt   = wplen   - wcnt;
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            wplen_nxt   = wplen      - wcnt;
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            wplen_nxt   = wplen;
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

assign tr_addrlsb_out = !(newCmd) ? addrlsb : tr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3 (
  input  wire            clk,
  input  wire            rst_n,
  // t
  output logic    [15:0] t_paddr,                                               // Address
  output logic           t_psel,                                                // Select
  output logic           t_penable,                                             // Enable
  output logic           t_pwrite,                                              // Write not read
  output logic    [31:0] t_pwdata,                                              // Write data
  output logic     [3:0] t_pstrb,                                               // Write strobes
  input  wire            t_pready,                                              // Ready
  input  wire     [31:0] t_prdata,                                              // Read data
  // f0
  input  wire            f0_activity,                                           // Upcoming activity indicator
  input  wire            f0_req,                                                // Flit transfer request
  input  wire            f0_sop,                                                // Start of packet indicator
  input  wire            f0_eop,                                                // End of packet indicator
  input  wire     [35:0] f0_flitdata,                                           // Flit data
  output logic           f0_ready,                                              // Flit transfer ready
  // f1
  input  wire            f1_activity,                                           // Upcoming activity indicator
  input  wire            f1_req,                                                // Flit transfer request
  input  wire            f1_sop,                                                // Start of packet indicator
  input  wire            f1_eop,                                                // End of packet indicator
  input  wire     [59:0] f1_flitdata,                                           // Flit data
  output logic           f1_ready,                                              // Flit transfer ready
  // r0
  output logic           r0_activity,                                           // Upcoming activity indicator
  output logic           r0_req,                                                // Flit transfer request
  output logic           r0_sop,                                                // Start of packet indicator
  output logic           r0_eop,                                                // End of packet indicator
  output logic    [33:0] r0_flitdata,                                           // Flit data
  input  wire            r0_ready,                                              // Flit transfer ready
  // r1
  output logic           r1_activity,                                           // Upcoming activity indicator
  output logic           r1_req,                                                // Flit transfer request
  output logic           r1_sop,                                                // Start of packet indicator
  output logic           r1_eop,                                                // End of packet indicator
  output logic    [23:0] r1_flitdata,                                           // Flit data
  input  wire            r1_ready                                               // Flit transfer ready
);

logic    [15:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic           wr_req;
logic           wr_ready;
logic           wr_last;
logic    [31:0] wr_data;
logic     [3:0] wr_strb;
logic           wc_buf_we;
logic    [71:0] wc_bus;
logic     [2:0] wc_sid;
logic     [2:0] wc_did;
logic     [1:0] wc_id;
logic    [31:0] wc_addr;
logic     [7:0] wc_len;
logic     [2:0] wc_rawsize;
logic     [2:0] wc_size;
logic     [1:0] wc_burst;
logic     [3:0] wc_qos;
logic     [2:0] wc_plen;
logic     [2:0] wc_prot;
logic           wcd_transinfo_en;
logic           wcd_transinfo_rdy;
logic           wf_req;
logic           wf_eop;
logic    [35:0] wf_flitdata;
logic           wf_ready;
logic    [23:0] ws_hdr;
logic           int_awvalid;
logic    [67:0] rds_hdr;
logic           rd_req;
logic           rd_ready;
logic           rd_last;
logic           rc_buf_we;
logic    [59:0] rc_bus;
logic     [2:0] rc_sid;
logic     [2:0] rc_did;
logic     [1:0] rc_id;
logic    [31:0] rc_addr;
logic     [2:0] rc_rawsize;
logic     [2:0] rc_size;
logic     [1:0] rc_burst;
logic     [3:0] rc_qos;
logic     [2:0] rc_plen;
logic     [2:0] rc_prot;
logic           rf_req;
logic           rf_eop;
logic    [33:0] rf_flitdata;
logic           rf_ready;
logic           rds_transinfo_we;
logic           rds_transinfo_rdy;
logic           int_arvalid;
logic    [11:0] wc_addr_unpack;
logic    [11:0] rc_addr_pack;
logic     [2:0] int_pprot;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           apbclk;
logic           apbclkAct;
logic           int_apbactivity;
logic           wcclk;
logic           wcclkAct;
wire            int_awactivity;
logic           wdclk;
logic           wdclkAct;
logic           int_wactivity;
logic           rcclk;
logic           rcclkAct;
logic           int_aractivity;
logic           rdclk;
logic           rdclkAct;
logic           rdclkEn;
logic           wrDone;
logic     [0:0] wr_cnt;
logic     [0:0] wr_cnt_nxt;
logic     [0:0] wr_cnt_en;
logic     [1:0] wr_state;
logic     [1:0] wr_state_nxt;
logic     [0:0] wr_state_en;
logic    [35:0] wc_buf [1:0];
logic     [1:0] wc_buf_en;
logic           int_pslverr;
logic     [0:0] rc_cnt;
logic     [0:0] rc_cnt_nxt;
logic     [0:0] rc_cnt_en;
logic           pslverr_w;
logic    [31:0] prdata;
logic     [1:0] rd_state;
logic     [1:0] rd_state_nxt;
logic     [0:0] rd_state_en;
logic    [59:0] rc_buf [0:0];
logic     [0:0] rc_buf_en;
logic           Narrow_Req;
logic     [1:0] apb_state;
logic     [1:0] apb_state_nxt;
logic     [0:0] apb_state_en;
logic     [0:0] apb_wrarb;
logic     [0:0] apb_wrarb_nxt;
logic     [0:0] apb_wrarb_en;
// ========================================================================//
// Parameter Declarations
// ========================================================================//
// ========================================================================//
// Process parameters and create local derived variables
// ========================================================================//
// ========================================================================//
// Define module I/O
// ========================================================================//
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Target Interface(s) (APB manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Egress APB Pipeline Component
usb4_tc_noc_apbtea3_epipe epipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(int_paddr),                                                        // i:16
  .src_psel(int_psel),                                                          // i:1
  .src_penable(int_penable),                                                    // i:1
  .src_pwrite(int_pwrite),                                                      // i:1
  .src_pwdata(int_pwdata),                                                      // i:32
  .src_pstrb(int_pstrb),                                                        // i:4
  .src_pready(int_pready),                                                      // o:1
  .src_prdata(int_prdata),                                                      // o:32
  .dst_paddr(t_paddr),                                                          // o:16
  .dst_psel(t_psel),                                                            // o:1
  .dst_penable(t_penable),                                                      // o:1
  .dst_pwrite(t_pwrite),                                                        // o:1
  .dst_pwdata(t_pwdata),                                                        // o:32
  .dst_pstrb(t_pstrb),                                                          // o:4
  .dst_pready(t_pready),                                                        // i:1
  .dst_prdata(t_prdata)                                                         // i:32
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea3_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f0_activity),                                                   // i:1
  .src_req(f0_req),                                                             // i:1
  .src_sop(f0_sop),                                                             // i:1
  .src_eop(f0_eop),                                                             // i:1
  .src_flitdata(f0_flitdata),                                                   // i:36
  .src_ready(f0_ready),                                                         // o:1
  .dst_activity(if0_activity),                                                  // o:1
  .dst_req(if0_req),                                                            // o:1
  .dst_sop(if0_sop),                                                            // o:1
  .dst_eop(if0_eop),                                                            // o:1
  .dst_flitdata(if0_flitdata),                                                  // o:36
  .dst_ready(if0_ready)                                                         // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea3_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f1_activity),                                                   // i:1
  .src_req(f1_req),                                                             // i:1
  .src_sop(f1_sop),                                                             // i:1
  .src_eop(f1_eop),                                                             // i:1
  .src_flitdata(f1_flitdata),                                                   // i:60
  .src_ready(f1_ready),                                                         // o:1
  .dst_activity(if1_activity),                                                  // o:1
  .dst_req(if1_req),                                                            // o:1
  .dst_sop(if1_sop),                                                            // o:1
  .dst_eop(if1_eop),                                                            // o:1
  .dst_flitdata(if1_flitdata),                                                  // o:60
  .dst_ready(if1_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea3_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir0_activity),                                                  // i:1
  .src_req(ir0_req),                                                            // i:1
  .src_sop(ir0_sop),                                                            // i:1
  .src_eop(ir0_eop),                                                            // i:1
  .src_flitdata(ir0_flitdata),                                                  // i:34
  .src_ready(ir0_ready),                                                        // o:1
  .dst_activity(r0_activity),                                                   // o:1
  .dst_req(r0_req),                                                             // o:1
  .dst_sop(r0_sop),                                                             // o:1
  .dst_eop(r0_eop),                                                             // o:1
  .dst_flitdata(r0_flitdata),                                                   // o:34
  .dst_ready(r0_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea3_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir1_activity),                                                  // i:1
  .src_req(ir1_req),                                                            // i:1
  .src_sop(ir1_sop),                                                            // i:1
  .src_eop(ir1_eop),                                                            // i:1
  .src_flitdata(ir1_flitdata),                                                  // i:24
  .src_ready(ir1_ready),                                                        // o:1
  .dst_activity(r1_activity),                                                   // o:1
  .dst_req(r1_req),                                                             // o:1
  .dst_sop(r1_sop),                                                             // o:1
  .dst_eop(r1_eop),                                                             // o:1
  .dst_flitdata(r1_flitdata),                                                   // o:24
  .dst_ready(r1_ready)                                                          // i:1
);
// =======================================================================
// Signal declarations
// =======================================================================
// Write Command + Data Sequencer Signals
// Write Command Signals
// Write Response Fields
// Read Data + Status fields
// Read Data + Status Flit Sequencer Signals
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea3_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign int_apbactivity = int_awactivity || int_aractivity;
usb4_tc_noc_apbtea3_apbcg apbcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_apbactivity),                                                      // i:1
  .clkOut(apbclk),                                                              // o:1
  .isActive(apbclkAct)                                                          // o:1
);
assign int_awactivity = if0_activity || if0_req || int_awvalid || ir1_req || wr_req;
usb4_tc_noc_apbtea3_wccg wccg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_awactivity),                                                       // i:1
  .clkOut(wcclk),                                                               // o:1
  .isActive(wcclkAct)                                                           // o:1
);
assign int_wactivity = if0_activity || if0_req || !wcd_transinfo_rdy || int_awvalid;
usb4_tc_noc_apbtea3_wdcg wdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_wactivity),                                                        // i:1
  .clkOut(wdclk),                                                               // o:1
  .isActive(wdclkAct)                                                           // o:1
);
assign ir1_activity = ir1_req;
assign int_aractivity = if1_activity || if1_req || ir0_req || rd_req;
usb4_tc_noc_apbtea3_f1cg f1cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_aractivity),                                                       // i:1
  .clkOut(rcclk),                                                               // o:1
  .isActive(rcclkAct)                                                           // o:1
);
assign ir0_activity = ir0_req;
assign rdclkEn = ir0_activity || if1_activity || if1_req || !rds_transinfo_rdy;
usb4_tc_noc_apbtea3_rdcg rdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(rdclkEn),                                                              // i:1
  .clkOut(rdclk),                                                               // o:1
  .isActive(rdclkAct)                                                           // o:1
);
// =======================================================================
// Write Processing
// =======================================================================
assign wrDone = wr_last && int_penable && int_pwrite && int_pready;
parameter S_WR_HDR = 2'd0;
parameter S_WR_DATA = 2'd1;
parameter S_WR_WAIT = 2'd2;
parameter S_WR_STS = 2'd3;
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign wc_bus[35:0] = wc_buf[0];
assign wc_bus[71:36] = ((wr_state == 2'b00) && (wr_cnt >= 1'd1)) ? if0_flitdata : wc_buf[1];
// Current Flit Count
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_cnt <= #1ps 1'd0;
  else if (wr_cnt_en)
    wr_cnt <= #1ps wr_cnt_nxt;
end

// Write State Machine State
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_state <= #1ps S_WR_HDR;
  else if (wr_state_en)
    wr_state <= #1ps wr_state_nxt;
end

// Write Command Packing Buffer
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      wc_buf[0] <= #1ps {36{1'b0}};
      wc_buf[1] <= #1ps {36{1'b0}};
    end
  else
    begin
      if (wc_buf_en[0])
        wc_buf[0] <= #1ps if0_flitdata;
      if (wc_buf_en[1])
        wc_buf[1] <= #1ps if0_flitdata;
    end
end

assign wc_buf_en = wc_buf_we << wr_cnt;
always_comb
begin
  // Defaults
  if0_ready    = 1'b0;
  ir1_req      = 1'b0;
  ir1_sop      = 1'b0;
  ir1_eop      = 1'b0;
  ir1_flitdata = {24{1'b0}};
  wr_cnt_nxt   = wr_cnt;
  wr_state_nxt = wr_state;
  wcd_transinfo_en = 1'b0;
  wf_req       = 1'b0;
  wf_eop       = 1'b0;
  wf_flitdata  = {36{1'b0}};
  // Write enables
  wc_buf_we    = 1'b0;
  wr_cnt_en    = 1'b0;
  wr_state_en  = 1'b0;
  int_awvalid   = 1'b0;
  case (wr_state)
    S_WR_HDR:
      begin
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_req)
          begin
            if0_ready    = 1'b1;
            // Header transmission is complete
            if (wr_cnt == 1'd1)
              begin
                int_awvalid = wcd_transinfo_rdy;
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wc_buf_we    = 1'b1;
                wcd_transinfo_en = 1'b1;
                wr_state_nxt = S_WR_DATA;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
                wc_buf_we  = 1'b1;
              end
          end
      end
   S_WR_DATA:
      begin
        wf_req      = if0_req;
        wf_eop      = if0_eop;
        wf_flitdata = if0_flitdata;
        if0_ready   = wf_ready;
        if (if0_req && wf_ready && if0_eop)
          begin
            wr_state_nxt = S_WR_WAIT;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_WAIT:
      begin
        if (wr_req && wr_ready && wr_last)
          begin
            wr_state_nxt = S_WR_STS;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_STS:
      begin
        ir1_req   = 1'b1;
        ir1_sop   = (wr_cnt == 1'd0);
        ir1_eop   = (wr_cnt == 1'd0);
        case(wr_cnt)
          1'd0: ir1_flitdata = ws_hdr[23:0];
          default: ir1_flitdata = {24{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_ready)
          begin
            // Header transmission is complete
            if (wr_cnt == 1'd0)
              begin
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wr_state_nxt = S_WR_HDR;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
              end
          end
      end
  endcase
end

 always_ff @(posedge wcclk) assert ( (frst_n===1'b0) || (int_awvalid == 1'b0) || (wc_burst != 2'b00) || ( {{(32-3){1'b0}},wc_plen} <= (32<<1) )) else $error("ERROR usb4_tc_noc_apbtea3 : %0t : Write data burst request is larger than TEA can handle. Write data burst size(wplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,wc_plen,(32<<1) );
usb4_tc_noc_apbtea3_wdunpack wdunpack (
  .clk(wdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .wtr_req(wcd_transinfo_en),                                                   // i:1
  .wtr_rdy(wcd_transinfo_rdy),                                                  // o:1
  .wtr_size(wc_size),                                                           // i:3
  .wtr_burst(wc_burst),                                                         // i:2
  .wtr_addrlsb(wc_addr[11:0]),                                                  // i:12
  .wtr_plen(wc_plen),                                                           // i:3
  .w_valid(wr_req),                                                             // o:1
  .w_data(wr_data),                                                             // o:32
  .w_strb(wr_strb),                                                             // o:4
  .w_last(wr_last),                                                             // o:1
  .w_ready(wr_ready),                                                           // i:1
  .f_req(wf_req),                                                               // i:1
  .f_eop(wf_eop),                                                               // i:1
  .f_flitdata(wf_flitdata),                                                     // i:36
  .f_ready(wf_ready),                                                           // o:1
  .wtr_addrlsb_out(wc_addr_unpack)                                              // o:12
);
// Write Command + Data Signal Unpacking
assign wc_sid = wc_bus[17:15];
assign wc_did = wc_bus[6:4];
assign wc_id = wc_bus[19:18];
assign wc_addr = wc_bus[54:23];
assign wc_qos = wc_bus[3:0];
assign wc_plen = wc_bus[22:20];
assign wc_prot = 3'd0;
assign wc_rawsize = wc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign wc_size = (wc_rawsize > 3'd2) ? 3'd2 : wc_rawsize;
assign wc_burst = wc_bus[59:58];
// =======================================================================
// Write Response Path Processing
// =======================================================================
// ============================================
// Write Response header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  ws_hdr            = {24{1'b0}};
  // Assign over the various fields
  ws_hdr[3:0]  = wc_qos;                                                        // loopback QoS from write command
  ws_hdr[6:4]  = wc_sid;                                                        // loopback SID from write command to DID
  ws_hdr[7]  = 1'b1;                                                            // SoT: not supporting fragmentation yet
  ws_hdr[8]  = 1'b1;                                                            // EoT: not supporting fragmentation yet
  ws_hdr[14:9]  = 6'd3;                                                         // Read command
  ws_hdr[17:15]  = wc_did;                                                      // loopback DID from wrtie command to SID
  ws_hdr[19:18]   = wc_id;
end

// declare the state parameters for read
parameter S_RC_HDR = 2'd0;
parameter S_RDS_WAIT = 2'd1;
parameter S_RDS_HDR = 2'd2;
parameter S_RDS_PLD = 2'd3;
assign int_pslverr = 1'd0;
// =======================================================================
// Read Processing
// =======================================================================
// Current Read Flit Count
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rc_cnt <= #1ps 1'd0;
  else if (rc_cnt_en)
    rc_cnt <= #1ps rc_cnt_nxt;
end

assign prdata = int_prdata;
assign pslverr_w = int_pslverr;
// Read State Machine State
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rd_state <= #1ps S_RC_HDR;
  else if (rd_state_en)
    rd_state <= #1ps rd_state_nxt;
end

// Read Command Packing Buffer
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rc_buf[0] <= #1ps {60{1'b0}};
    end
  else
    begin
      if (rc_buf_en[0])
        rc_buf[0] <= #1ps if1_flitdata;
    end
end

assign rc_buf_en = rc_buf_we << rc_cnt;
// ============================================
// Read Data + Status flit sequencer
// ============================================
always_comb
begin
  // Defaults
  rd_state_nxt  = rd_state;
  rc_cnt_nxt    = rc_cnt;
  ir0_req       = 1'b0;
  ir0_sop       = 1'b0;
  ir0_eop       = 1'b0;
  ir0_flitdata  = {34{1'b0}};
  rds_transinfo_we = 1'b0;
  if1_ready     = 1'b0;
  rf_ready      = 1'b0;
  // Write enables
  rd_state_en   = 1'b0;
  rc_cnt_en     = 1'b0;
  rc_buf_we     = 1'b0;
  int_arvalid  = 1'b0;
  case (rd_state)
    S_RC_HDR:
      begin
        if1_ready    = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if1_req)
          begin
            // Header transmission is complete
            if (rc_cnt == 1'd0)
              begin
                int_arvalid  = 1'b1;
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rc_buf_we    = 1'b1;
                rds_transinfo_we = 1'b1;
                rd_state_nxt = S_RDS_WAIT;
                rd_state_en   = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                rc_buf_we    = 1'b1;
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
   S_RDS_WAIT:
   begin
    if (int_pready && int_penable && !int_pwrite)
    begin
        rd_state_nxt = S_RDS_HDR;
        rd_state_en  = 1'b1;
    end
   end
   S_RDS_HDR:
      begin
        ir0_req   = 1'd1;
        ir0_sop   = (rc_cnt == 1'd0);
        case(rc_cnt)
          1'd0: ir0_flitdata = rds_hdr[33:0];
          1'd1: ir0_flitdata = rds_hdr[67:34];
          default: ir0_flitdata = {34{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir0_req && ir0_ready)
          begin
            // Complete header is done
            if (rc_cnt == 1'd1)
              begin
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rd_state_nxt = S_RDS_PLD;
                rd_state_en   = 1'b1;
              end
            else
              begin
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
    S_RDS_PLD:
      begin
        ir0_req       = rf_req;
        ir0_eop       = rf_eop;
        ir0_flitdata  = rf_flitdata;
        rf_ready      = ir0_ready;
        if (rf_req && rf_eop && ir0_ready)
          begin
            rd_state_nxt = S_RC_HDR;
            rd_state_en   = 1'b1;
          end
      end
  endcase
end

always_ff @(posedge rcclk) assert ( (frst_n===1'b0) || (int_arvalid == 1'b0) || (rc_burst != 2'b00) || ({{(32-3){1'b0}},rc_plen} <= (32<<1) ) ) else $error("ERROR usb4_tc_noc_apbtea3 : %0t : Read data burst request is larger than TEA can handle. Read data burst size(rplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,rc_plen,(32<<1) );
usb4_tc_noc_apbtea3_rdpack rdpack (
  .clk(rdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .tr_req(rds_transinfo_we),                                                    // i:1
  .tr_rdy(rds_transinfo_rdy),                                                   // o:1
  .tr_size(rc_size),                                                            // i:3
  .tr_burst(rc_burst),                                                          // i:2
  .tr_addrlsb(rc_addr[11:0]),                                                   // i:12
  .tr_plen(rc_plen),                                                            // i:3
  .r_req(rd_req),                                                               // o:1
  .r_last(rd_last),                                                             // o:1
  .r_data(prdata),                                                              // i:32
  .r_slverr(pslverr_w),                                                         // i:1
  .r_ready(rd_ready),                                                           // i:1
  .f_req(rf_req),                                                               // o:1
  .f_eop(rf_eop),                                                               // o:1
  .f_flitdata(rf_flitdata),                                                     // o:34
  .f_ready(rf_ready),                                                           // i:1
  .tr_addrlsb_out(rc_addr_pack)                                                 // o:12
);
// Create incoming rc bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rc_bus[59:0] = (rd_state == S_RC_HDR) ? if1_flitdata : rc_buf[0];
// assign rc.bus = {$rcBusStr};
// Read Command Signal Unpacking
assign rc_sid = rc_bus[17:15];
assign rc_did = rc_bus[6:4];
assign rc_id = rc_bus[19:18];
assign rc_addr = rc_bus[54:23];
assign rc_qos = rc_bus[3:0];
assign rc_plen = rc_bus[22:20];
assign rc_prot = 3'd0;
assign rc_rawsize = rc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign rc_size = Narrow_Req ? ((rc_rawsize < 3'd2) ? rc_rawsize : 3'd2) : ((rc_rawsize > 3'd2) ? 3'd2 : rc_rawsize);
assign rc_burst = rc_bus[59:58];
assign Narrow_Req = rc_rawsize < 3'd2;
// ============================================
// Read Data + Status Header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  rds_hdr            = {68{1'b0}};
  // Assign over the various fields
  rds_hdr[3:0]  = rc_qos;                                                       // loopback QoS from write command
  rds_hdr[6:4]  = rc_sid;                                                       // loopback SID from write command to DID
  rds_hdr[7]  = 1'b1;                                                           // SoT: not supporting fragmentation yet
  rds_hdr[8]  = 1'b1;                                                           // EoT: not supporting fragmentation yet
  rds_hdr[14:9]  = 6'd1;                                                        // Read data / status
  rds_hdr[17:15]  = rc_did;                                                     // loopback DID from wrtie command to SID
  rds_hdr[19:18]   = rc_id;
  rds_hdr[22:20] = rc_plen;
  rds_hdr[30:23]  = (rc_burst==2'd2) ? 8'(rc_addr[11:0] >> rc_size) : rc_addr[7:0];
  rds_hdr[33:31]  = rc_size;
  rds_hdr[35:34] = rc_burst;
end

// Arbitrate between read and write state machines for use of APB interface
parameter S_PSEL = 2'd0;
parameter S_PWEN = 2'd1;
parameter S_PREN = 2'd2;
parameter S_PRDATA = 2'd3;
// APB State Machine State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_state <= #1ps S_PSEL;
  else if (apb_state_en)
    apb_state <= #1ps apb_state_nxt;
end

// Read / Write Arbiter State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_wrarb <= #1ps 1'd0;
  else if (apb_wrarb_en)
    apb_wrarb <= #1ps apb_wrarb_nxt;
end

// For multiple targets and when both rd and wr are active
always_comb
begin
  int_psel      = 1'b0;
  int_pwrite    = 1'b0;
  int_penable   = 1'b0;
  int_paddr     = {16{1'b0}};
  int_pwdata    = {32{1'b0}};
  int_pstrb     = {4{1'b0}};
  int_pprot     = 3'd0;
  apb_state_nxt = apb_state;
  apb_state_en  = 1'b0;
  apb_wrarb_nxt = apb_wrarb;
  apb_wrarb_en  = 1'b0;
  wr_ready      = 1'b0;
  rd_ready      = 1'b0;
  case (apb_state)
    S_PSEL:
      begin
        if (wr_req && (!rd_req || apb_wrarb))
          begin
            int_psel      = 1'b1;
            int_paddr     = {wc_addr[15:12],wc_addr_unpack};
            int_pwrite    = 1'b1;
            int_pwdata    = wr_data;
            int_pstrb     = wr_strb;
            int_pprot     = wc_prot;
            apb_state_nxt = S_PWEN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b0;
            apb_wrarb_en  = 1'b1;
          end
        else if (rd_req)
          begin
            int_psel      = 1'b1;
            int_paddr     = {rc_addr[15:12],rc_addr_pack};
            int_pprot     = rc_prot;
            apb_state_nxt = S_PREN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b1;
            apb_wrarb_en  = 1'b1;
          end
      end
    S_PWEN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
        int_pwrite  = 1'b1;
        int_paddr   = {wc_addr[15:12],wc_addr_unpack};
        int_pwdata  = wr_data;
        int_pstrb   = wr_strb;
        int_pprot   = wc_prot;
        if (int_pready)
          begin
            wr_ready   = 1'b1;
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
          end
      end
    S_PREN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
            int_paddr     = {rc_addr[15:12],rc_addr_pack};
        int_pprot   = rc_prot;
        if (int_pready)
          begin
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
            rd_ready   = 1'b1;
          end
      end
    // S_PRDATA:
    // begin
    // apb.state.nxt = S_PSEL;
    // apb.state.en  = 1'b1;
    // end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_epipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire     [15:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  // dst
  output logic    [15:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata                                             // Read data
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea3_epipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_epipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea3_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea3_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea3_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea3_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_apbcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_wccg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_wdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_f1cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_rdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_wdunpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wtr_req,
  output logic           wtr_rdy,
  input  wire      [2:0] wtr_size,                                              // Transfer size per data phase
  input  wire      [1:0] wtr_burst,                                             // Burst addressing mode
  input  wire     [11:0] wtr_addrlsb,                                           // 12 LSBs of address
  input  wire      [2:0] wtr_plen,                                              // Packet length in bytes
  output logic           w_valid,
  output logic    [31:0] w_data,
  output logic     [3:0] w_strb,
  output logic           w_last,
  input  wire            w_ready,
  input  wire            f_req,
  input  wire            f_eop,
  input  wire     [35:0] f_flitdata,
  output logic           f_ready,
  output logic    [11:0] wtr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [2:0] sizeCnvDiv;
logic     [4:0] firstCnt2Wrap;
logic     [7:0] wtr_mask;
logic     [7:0] wtr_mis;
logic    [10:0] firstXferCnt;
logic    [10:0] xferCnt;
logic    [10:0] xferCnt_nxt;
logic     [0:0] xferCnt_en;
logic    [10:0] useXferCnt;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic    [31:0] muxed_w_data;
logic     [3:0] muxed_w_strb;
logic           flitDone;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic     [0:0] haveFlit;
logic     [0:0] haveFlit_nxt;
logic     [0:0] haveFlit_en;
logic    [35:0] flitData;
logic    [35:0] flitData_nxt;
logic     [0:0] flitData_en;
logic           flitValid;
logic    [11:0] lower_baddr;
logic    [11:0] upper_baddr;
logic    [11:0] lower_addr;
logic    [11:0] upper_addr;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
logic    [11:0] saddr;
logic     [2:0] splen;
// Extracted from packet header
// APB W Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},wtr_plen} - 1'b1;                                    // We only care about 8 bits of address for our word indexing
assign wrapToAddr = wtr_addrlsb[7:0] & ~bamask;                                 // This is the address offset we wrap to
assign wrapIndex = wtr_addrlsb >> wtr_size;
assign sizeCnvDiv = wtr_plen >> wtr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign wtr_mask = (8'b1<<wtr_size) - 1'b1;
assign wtr_mis = wtr_addrlsb[7:0] & wtr_mask;
assign firstXferCnt = (wtr_burst!=2'd1) ? 11'(wtr_plen>>wtr_size) : 11'((16'(wtr_plen)+wtr_mask+wtr_mis)>>wtr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    xferCnt <= #1ps 11'd0;
  else if (xferCnt_en)
    xferCnt <= #1ps xferCnt_nxt;
end

assign useXferCnt = xferCnt;
always_comb
begin
  xferCnt_nxt = xferCnt;
  xferCnt_en  = 1'b0;
  if( newCmd )
    begin
      xferCnt_nxt = firstXferCnt;
      xferCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      xferCnt_nxt = useXferCnt - 1'd1;
      xferCnt_en  = 1'b1;
    end
end

assign wtr_rdy = ~trInPkt;
assign newCmd = wtr_req && wtr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = w_valid && w_ready;
assign f_ready = ~haveFlit || flitDone;
assign w_valid = flitValid;
assign w_last = w_valid && useXferCnt==11'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps wtr_burst;
end

assign use_tr_burst = held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps wtr_size;
end

assign use_tr_size = held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( busWriteValid && w_last )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> wtr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (wtr_addrlsb[7:0] & 8'd3) >> wtr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( w_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone;
assign muxed_w_data[7:0] = flitData[7:0];
assign muxed_w_strb[3:0] = flitData[35:32];
assign muxed_w_data[15:8] = flitData[15:8];
assign muxed_w_data[23:16] = flitData[23:16];
assign muxed_w_data[31:24] = flitData[31:24];
assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    haveFlit <= #1ps 1'd0;
  else if (haveFlit_en)
    haveFlit <= #1ps haveFlit_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitData <= #1ps {36{1'b0}};
  else if (flitData_en)
    flitData <= #1ps flitData_nxt;
end

assign flitValid = haveFlit;
always_comb
begin
  haveFlit_nxt   = haveFlit;
  haveFlit_en    = 1'b0;
  flitData_nxt   = flitData;
  flitData_en    = 1'b0;
  if( flitWriteValid )
    begin
      haveFlit_nxt   = 1'b1;
      haveFlit_en    = 1'b1;
      flitData_en    = 1'b1;
      flitData_nxt   = f_flitdata;
    end
  else if( flitDone )
    begin
      haveFlit_nxt   = 1'b0;
      haveFlit_en    = 1'b1;
    end
end

assign w_data[7:0] = (w_valid && wrMask[0]) ? muxed_w_data[7:0] : 8'd0;
assign w_data[15:8] = (w_valid && wrMask[1]) ? muxed_w_data[15:8] : 8'd0;
assign w_data[23:16] = (w_valid && wrMask[2]) ? muxed_w_data[23:16] : 8'd0;
assign w_data[31:24] = (w_valid && wrMask[3]) ? muxed_w_data[31:24] : 8'd0;
assign w_strb = w_valid ? muxed_w_strb & wrMask : 4'd0;
assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  addrlsb_nxt   = addrlsb;
  // Write enables
  addrlsb_en    = 1'b0;
  if (newCmd)
    begin
      addrlsb_nxt = wtr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred from packing FIFO
  else if (busWriteValid)
    begin
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps wtr_addrlsb;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps wtr_plen;
end

assign wtr_addrlsb_out = !(newCmd) ? addrlsb : wtr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea3_rdpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            tr_req,
  output logic           tr_rdy,
  input  wire      [2:0] tr_size,
  input  wire      [1:0] tr_burst,
  input  wire     [11:0] tr_addrlsb,
  input  wire      [2:0] tr_plen,
  output logic           r_req,
  output logic           r_last,
  input  wire     [31:0] r_data,
  input  wire            r_slverr,
  input  wire            r_ready,
  output logic           f_req,
  output logic           f_eop,
  output logic    [33:0] f_flitdata,
  input  wire            f_ready,
  output logic    [11:0] tr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [4:0] firstCnt2Wrap;
logic     [2:0] sizeCnvDiv;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [0:0] heldFlitDone;
logic     [0:0] heldEop;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isNarrow;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic           flitDone;
logic           useBusWdCnt;
logic    [33:0] flitWd;
logic    [33:0] flitWd_nxt;
logic     [0:0] flitWd_en;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] lower_baddr;                                                    // Lower burst address
logic    [11:0] upper_baddr;                                                    // Upper burst address
logic    [11:0] lower_addr;                                                     // Lower element address
logic    [11:0] upper_addr;                                                     // Upper element address
logic    [11:0] esize_minus_first_offset;
logic    [11:0] first_offset;
logic     [2:0] raw_wcnt;
logic     [2:0] wcnt;
logic    [11:0] saddr;
logic     [2:0] wplen;
logic     [2:0] wplen_nxt;
logic     [0:0] wplen_en;
logic     [2:0] splen;
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
// Extracted from AXI AW Channel
// APB R Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},tr_plen} - 1'b1;                                     // We only care about 8 bits of address for our word indexing
assign wrapToAddr = tr_addrlsb[7:0] & ~bamask;                                  // This is the address offset we wrap to
assign wrapIndex = tr_addrlsb >> tr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign sizeCnvDiv = tr_plen >> tr_size;
assign tr_rdy = ~trInPkt;
assign f_flitdata = flitWd;
assign f_req = heldFlitDone;
assign f_eop = heldEop;
assign r_req = trInPkt_nxt && (!heldFlitDone || flitWriteValid);
assign newCmd = tr_req && tr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = r_ready && r_req;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldFlitDone <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldFlitDone <= #1ps flitDone;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldEop <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldEop <= #1ps flitDone && r_last;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps tr_burst;
end

assign use_tr_burst = (newCmd) ? tr_burst : held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps tr_size;
end

assign use_tr_size = (newCmd) ? tr_size : held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isNarrow = use_tr_size<3'd2;
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( flitWriteValid && f_eop )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> tr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = (newCmd) ? subBusWdCntWrap_nxt : subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = newCmd ? firstCnt2Wrap : cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (tr_addrlsb[7:0] & 8'd3) >> tr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = (newCmd) ? firstSubBusWdCnt[1:0] : subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( r_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone || (isNarrow && busWriteValid);
assign useBusWdCnt = 1'b0;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitWd <= #1ps {34{1'b0}};
  else if (flitWd_en)
    flitWd <= #1ps flitWd_nxt;
end

assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_comb
begin
  // First, assign the bus word to every possible flit word slot
  flitWd_nxt = flitWriteValid ? {34{1'b0}} : flitWd;
  // Start out with nothing enabled
  flitWd_en = flitWriteValid ? 1'b1 : 1'b0;
  // Now enable any bytes that are being written this cycle
  if( busWriteValid )
    begin
      if( useBusWdCnt == 1'd0 )
        begin
          if( wrMask[0] )
            begin
              flitWd_nxt[7:0] = r_data[7:0];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[1] )
            begin
              flitWd_nxt[15:8] = r_data[15:8];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[2] )
            begin
              flitWd_nxt[23:16] = r_data[23:16];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[3] )
            begin
              flitWd_nxt[31:24] = r_data[31:24];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
        end
    end
end

assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
assign esize_minus_first_offset = esize - first_offset;
assign first_offset = addrlsb & amask;
assign raw_wcnt = (held_tr_burst == 2'd1) ? esize_minus_first_offset[2:0] : esize[2:0];
assign wcnt = (raw_wcnt > wplen) ? wplen : raw_wcnt;
assign r_last = (wcnt >= wplen);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps tr_addrlsb;
end

// Write remaining packet length and address LSB tracking flops
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    wplen <= #1ps 3'd0;
  else if (wplen_en)
    wplen <= #1ps wplen_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps tr_plen;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  wplen_nxt   = wplen;
  addrlsb_nxt = addrlsb;
  wplen_en    = 1'b0;
  addrlsb_en  = 1'b0;
  if (tr_req && tr_rdy)
    begin
      wplen_nxt   = tr_plen;
      wplen_en    = 1'b1;
      addrlsb_nxt = tr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred to packing FIFO
  else if (busWriteValid)
    begin
      wplen_en    = 1'b1;
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            wplen_nxt   = wplen - wcnt;
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            wplen_nxt   = wplen   - wcnt;
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            wplen_nxt   = wplen      - wcnt;
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            wplen_nxt   = wplen;
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

assign tr_addrlsb_out = !(newCmd) ? addrlsb : tr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4 (
  input  wire            clk,
  input  wire            rst_n,
  // t
  output logic    [17:0] t_paddr,                                               // Address
  output logic           t_psel,                                                // Select
  output logic           t_penable,                                             // Enable
  output logic           t_pwrite,                                              // Write not read
  output logic    [31:0] t_pwdata,                                              // Write data
  output logic     [3:0] t_pstrb,                                               // Write strobes
  input  wire            t_pready,                                              // Ready
  input  wire     [31:0] t_prdata,                                              // Read data
  input  wire            t_pslverr,                                             // Slave error
  // f0
  input  wire            f0_activity,                                           // Upcoming activity indicator
  input  wire            f0_req,                                                // Flit transfer request
  input  wire            f0_sop,                                                // Start of packet indicator
  input  wire            f0_eop,                                                // End of packet indicator
  input  wire     [35:0] f0_flitdata,                                           // Flit data
  output logic           f0_ready,                                              // Flit transfer ready
  // f1
  input  wire            f1_activity,                                           // Upcoming activity indicator
  input  wire            f1_req,                                                // Flit transfer request
  input  wire            f1_sop,                                                // Start of packet indicator
  input  wire            f1_eop,                                                // End of packet indicator
  input  wire     [59:0] f1_flitdata,                                           // Flit data
  output logic           f1_ready,                                              // Flit transfer ready
  // r0
  output logic           r0_activity,                                           // Upcoming activity indicator
  output logic           r0_req,                                                // Flit transfer request
  output logic           r0_sop,                                                // Start of packet indicator
  output logic           r0_eop,                                                // End of packet indicator
  output logic    [33:0] r0_flitdata,                                           // Flit data
  input  wire            r0_ready,                                              // Flit transfer ready
  // r1
  output logic           r1_activity,                                           // Upcoming activity indicator
  output logic           r1_req,                                                // Flit transfer request
  output logic           r1_sop,                                                // Start of packet indicator
  output logic           r1_eop,                                                // End of packet indicator
  output logic    [23:0] r1_flitdata,                                           // Flit data
  input  wire            r1_ready                                               // Flit transfer ready
);

logic    [17:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           int_pslverr;                                                    // Slave error
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic           wr_req;
logic           wr_ready;
logic           wr_last;
logic    [31:0] wr_data;
logic     [3:0] wr_strb;
logic           wc_buf_we;
logic    [71:0] wc_bus;
logic     [2:0] wc_sid;
logic     [2:0] wc_did;
logic     [1:0] wc_id;
logic    [31:0] wc_addr;
logic     [7:0] wc_len;
logic     [2:0] wc_rawsize;
logic     [2:0] wc_size;
logic     [1:0] wc_burst;
logic     [3:0] wc_qos;
logic     [2:0] wc_plen;
logic     [2:0] wc_prot;
logic           wcd_transinfo_en;
logic           wcd_transinfo_rdy;
logic           wf_req;
logic           wf_eop;
logic    [35:0] wf_flitdata;
logic           wf_ready;
logic    [23:0] ws_hdr;
logic           int_awvalid;
logic    [67:0] rds_hdr;
logic           rd_req;
logic           rd_ready;
logic           rd_last;
logic           rc_buf_we;
logic    [59:0] rc_bus;
logic     [2:0] rc_sid;
logic     [2:0] rc_did;
logic     [1:0] rc_id;
logic    [31:0] rc_addr;
logic     [2:0] rc_rawsize;
logic     [2:0] rc_size;
logic     [1:0] rc_burst;
logic     [3:0] rc_qos;
logic     [2:0] rc_plen;
logic     [2:0] rc_prot;
logic           rf_req;
logic           rf_eop;
logic    [33:0] rf_flitdata;
logic           rf_ready;
logic           rds_transinfo_we;
logic           rds_transinfo_rdy;
logic           int_arvalid;
logic     [3:0] pslverrWr_4bit;
logic     [3:0] pslverrRd_4bit;
logic    [11:0] wc_addr_unpack;
logic    [11:0] rc_addr_pack;
logic     [2:0] int_pprot;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           apbclk;
logic           apbclkAct;
logic           int_apbactivity;
logic           wcclk;
logic           wcclkAct;
wire            int_awactivity;
logic           wdclk;
logic           wdclkAct;
logic           int_wactivity;
logic           rcclk;
logic           rcclkAct;
logic           int_aractivity;
logic           rdclk;
logic           rdclkAct;
logic           rdclkEn;
logic           wrDone;
logic     [0:0] wr_cnt;
logic     [0:0] wr_cnt_nxt;
logic     [0:0] wr_cnt_en;
logic     [1:0] wr_state;
logic     [1:0] wr_state_nxt;
logic     [0:0] wr_state_en;
logic    [35:0] wc_buf [1:0];
logic     [1:0] wc_buf_en;
logic           setWrError;
logic           clrWrError;
logic     [0:0] pslverrWr_latch;
logic     [0:0] pslverrWr_latch_nxt;
logic           setRdError;
logic           clrRdError;
logic     [0:0] pslverrRd_latch;
logic     [0:0] pslverrRd_latch_nxt;
logic     [0:0] rc_cnt;
logic     [0:0] rc_cnt_nxt;
logic     [0:0] rc_cnt_en;
logic           pslverr_w;
logic    [31:0] prdata;
logic     [1:0] rd_state;
logic     [1:0] rd_state_nxt;
logic     [0:0] rd_state_en;
logic    [59:0] rc_buf [0:0];
logic     [0:0] rc_buf_en;
logic           Narrow_Req;
logic     [1:0] apb_state;
logic     [1:0] apb_state_nxt;
logic     [0:0] apb_state_en;
logic     [0:0] apb_wrarb;
logic     [0:0] apb_wrarb_nxt;
logic     [0:0] apb_wrarb_en;
// ========================================================================//
// Parameter Declarations
// ========================================================================//
// ========================================================================//
// Process parameters and create local derived variables
// ========================================================================//
// ========================================================================//
// Define module I/O
// ========================================================================//
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Target Interface(s) (APB manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Egress APB Pipeline Component
usb4_tc_noc_apbtea4_epipe epipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(int_paddr),                                                        // i:18
  .src_psel(int_psel),                                                          // i:1
  .src_penable(int_penable),                                                    // i:1
  .src_pwrite(int_pwrite),                                                      // i:1
  .src_pwdata(int_pwdata),                                                      // i:32
  .src_pstrb(int_pstrb),                                                        // i:4
  .src_pready(int_pready),                                                      // o:1
  .src_prdata(int_prdata),                                                      // o:32
  .src_pslverr(int_pslverr),                                                    // o:1
  .dst_paddr(t_paddr),                                                          // o:18
  .dst_psel(t_psel),                                                            // o:1
  .dst_penable(t_penable),                                                      // o:1
  .dst_pwrite(t_pwrite),                                                        // o:1
  .dst_pwdata(t_pwdata),                                                        // o:32
  .dst_pstrb(t_pstrb),                                                          // o:4
  .dst_pready(t_pready),                                                        // i:1
  .dst_prdata(t_prdata),                                                        // i:32
  .dst_pslverr(t_pslverr)                                                       // i:1
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea4_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f0_activity),                                                   // i:1
  .src_req(f0_req),                                                             // i:1
  .src_sop(f0_sop),                                                             // i:1
  .src_eop(f0_eop),                                                             // i:1
  .src_flitdata(f0_flitdata),                                                   // i:36
  .src_ready(f0_ready),                                                         // o:1
  .dst_activity(if0_activity),                                                  // o:1
  .dst_req(if0_req),                                                            // o:1
  .dst_sop(if0_sop),                                                            // o:1
  .dst_eop(if0_eop),                                                            // o:1
  .dst_flitdata(if0_flitdata),                                                  // o:36
  .dst_ready(if0_ready)                                                         // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea4_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f1_activity),                                                   // i:1
  .src_req(f1_req),                                                             // i:1
  .src_sop(f1_sop),                                                             // i:1
  .src_eop(f1_eop),                                                             // i:1
  .src_flitdata(f1_flitdata),                                                   // i:60
  .src_ready(f1_ready),                                                         // o:1
  .dst_activity(if1_activity),                                                  // o:1
  .dst_req(if1_req),                                                            // o:1
  .dst_sop(if1_sop),                                                            // o:1
  .dst_eop(if1_eop),                                                            // o:1
  .dst_flitdata(if1_flitdata),                                                  // o:60
  .dst_ready(if1_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea4_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir0_activity),                                                  // i:1
  .src_req(ir0_req),                                                            // i:1
  .src_sop(ir0_sop),                                                            // i:1
  .src_eop(ir0_eop),                                                            // i:1
  .src_flitdata(ir0_flitdata),                                                  // i:34
  .src_ready(ir0_ready),                                                        // o:1
  .dst_activity(r0_activity),                                                   // o:1
  .dst_req(r0_req),                                                             // o:1
  .dst_sop(r0_sop),                                                             // o:1
  .dst_eop(r0_eop),                                                             // o:1
  .dst_flitdata(r0_flitdata),                                                   // o:34
  .dst_ready(r0_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea4_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir1_activity),                                                  // i:1
  .src_req(ir1_req),                                                            // i:1
  .src_sop(ir1_sop),                                                            // i:1
  .src_eop(ir1_eop),                                                            // i:1
  .src_flitdata(ir1_flitdata),                                                  // i:24
  .src_ready(ir1_ready),                                                        // o:1
  .dst_activity(r1_activity),                                                   // o:1
  .dst_req(r1_req),                                                             // o:1
  .dst_sop(r1_sop),                                                             // o:1
  .dst_eop(r1_eop),                                                             // o:1
  .dst_flitdata(r1_flitdata),                                                   // o:24
  .dst_ready(r1_ready)                                                          // i:1
);
// =======================================================================
// Signal declarations
// =======================================================================
// Write Command + Data Sequencer Signals
// Write Command Signals
// Write Response Fields
// Read Data + Status fields
// Read Data + Status Flit Sequencer Signals
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea4_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign int_apbactivity = int_awactivity || int_aractivity;
usb4_tc_noc_apbtea4_apbcg apbcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_apbactivity),                                                      // i:1
  .clkOut(apbclk),                                                              // o:1
  .isActive(apbclkAct)                                                          // o:1
);
assign int_awactivity = if0_activity || if0_req || int_awvalid || ir1_req || wr_req;
usb4_tc_noc_apbtea4_wccg wccg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_awactivity),                                                       // i:1
  .clkOut(wcclk),                                                               // o:1
  .isActive(wcclkAct)                                                           // o:1
);
assign int_wactivity = if0_activity || if0_req || !wcd_transinfo_rdy || int_awvalid;
usb4_tc_noc_apbtea4_wdcg wdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_wactivity),                                                        // i:1
  .clkOut(wdclk),                                                               // o:1
  .isActive(wdclkAct)                                                           // o:1
);
assign ir1_activity = ir1_req;
assign int_aractivity = if1_activity || if1_req || ir0_req || rd_req;
usb4_tc_noc_apbtea4_f1cg f1cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_aractivity),                                                       // i:1
  .clkOut(rcclk),                                                               // o:1
  .isActive(rcclkAct)                                                           // o:1
);
assign ir0_activity = ir0_req;
assign rdclkEn = ir0_activity || if1_activity || if1_req || !rds_transinfo_rdy;
usb4_tc_noc_apbtea4_rdcg rdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(rdclkEn),                                                              // i:1
  .clkOut(rdclk),                                                               // o:1
  .isActive(rdclkAct)                                                           // o:1
);
// =======================================================================
// Write Processing
// =======================================================================
assign wrDone = wr_last && int_penable && int_pwrite && int_pready;
parameter S_WR_HDR = 2'd0;
parameter S_WR_DATA = 2'd1;
parameter S_WR_WAIT = 2'd2;
parameter S_WR_STS = 2'd3;
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign wc_bus[35:0] = wc_buf[0];
assign wc_bus[71:36] = ((wr_state == 2'b00) && (wr_cnt >= 1'd1)) ? if0_flitdata : wc_buf[1];
// Current Flit Count
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_cnt <= #1ps 1'd0;
  else if (wr_cnt_en)
    wr_cnt <= #1ps wr_cnt_nxt;
end

// Write State Machine State
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_state <= #1ps S_WR_HDR;
  else if (wr_state_en)
    wr_state <= #1ps wr_state_nxt;
end

// Write Command Packing Buffer
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      wc_buf[0] <= #1ps {36{1'b0}};
      wc_buf[1] <= #1ps {36{1'b0}};
    end
  else
    begin
      if (wc_buf_en[0])
        wc_buf[0] <= #1ps if0_flitdata;
      if (wc_buf_en[1])
        wc_buf[1] <= #1ps if0_flitdata;
    end
end

assign wc_buf_en = wc_buf_we << wr_cnt;
always_comb
begin
  // Defaults
  if0_ready    = 1'b0;
  ir1_req      = 1'b0;
  ir1_sop      = 1'b0;
  ir1_eop      = 1'b0;
  ir1_flitdata = {24{1'b0}};
  wr_cnt_nxt   = wr_cnt;
  wr_state_nxt = wr_state;
  wcd_transinfo_en = 1'b0;
  wf_req       = 1'b0;
  wf_eop       = 1'b0;
  wf_flitdata  = {36{1'b0}};
  // Write enables
  wc_buf_we    = 1'b0;
  wr_cnt_en    = 1'b0;
  wr_state_en  = 1'b0;
  int_awvalid   = 1'b0;
  case (wr_state)
    S_WR_HDR:
      begin
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_req)
          begin
            if0_ready    = 1'b1;
            // Header transmission is complete
            if (wr_cnt == 1'd1)
              begin
                int_awvalid = wcd_transinfo_rdy;
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wc_buf_we    = 1'b1;
                wcd_transinfo_en = 1'b1;
                wr_state_nxt = S_WR_DATA;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
                wc_buf_we  = 1'b1;
              end
          end
      end
   S_WR_DATA:
      begin
        wf_req      = if0_req;
        wf_eop      = if0_eop;
        wf_flitdata = if0_flitdata;
        if0_ready   = wf_ready;
        if (if0_req && wf_ready && if0_eop)
          begin
            wr_state_nxt = S_WR_WAIT;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_WAIT:
      begin
        if (wr_req && wr_ready && wr_last)
          begin
            wr_state_nxt = S_WR_STS;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_STS:
      begin
        ir1_req   = 1'b1;
        ir1_sop   = (wr_cnt == 1'd0);
        ir1_eop   = (wr_cnt == 1'd0);
        case(wr_cnt)
          1'd0: ir1_flitdata = ws_hdr[23:0];
          default: ir1_flitdata = {24{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_ready)
          begin
            // Header transmission is complete
            if (wr_cnt == 1'd0)
              begin
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wr_state_nxt = S_WR_HDR;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
              end
          end
      end
  endcase
end

 always_ff @(posedge wcclk) assert ( (frst_n===1'b0) || (int_awvalid == 1'b0) || (wc_burst != 2'b00) || ( {{(32-3){1'b0}},wc_plen} <= (32<<1) )) else $error("ERROR usb4_tc_noc_apbtea4 : %0t : Write data burst request is larger than TEA can handle. Write data burst size(wplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,wc_plen,(32<<1) );
usb4_tc_noc_apbtea4_wdunpack wdunpack (
  .clk(wdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .wtr_req(wcd_transinfo_en),                                                   // i:1
  .wtr_rdy(wcd_transinfo_rdy),                                                  // o:1
  .wtr_size(wc_size),                                                           // i:3
  .wtr_burst(wc_burst),                                                         // i:2
  .wtr_addrlsb(wc_addr[11:0]),                                                  // i:12
  .wtr_plen(wc_plen),                                                           // i:3
  .w_valid(wr_req),                                                             // o:1
  .w_data(wr_data),                                                             // o:32
  .w_strb(wr_strb),                                                             // o:4
  .w_last(wr_last),                                                             // o:1
  .w_ready(wr_ready),                                                           // i:1
  .f_req(wf_req),                                                               // i:1
  .f_eop(wf_eop),                                                               // i:1
  .f_flitdata(wf_flitdata),                                                     // i:36
  .f_ready(wf_ready),                                                           // o:1
  .wtr_addrlsb_out(wc_addr_unpack)                                              // o:12
);
// Write Command + Data Signal Unpacking
assign wc_sid = wc_bus[17:15];
assign wc_did = wc_bus[6:4];
assign wc_id = wc_bus[19:18];
assign wc_addr = wc_bus[54:23];
assign wc_qos = wc_bus[3:0];
assign wc_plen = wc_bus[22:20];
assign wc_prot = 3'd0;
assign wc_rawsize = wc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign wc_size = (wc_rawsize > 3'd2) ? 3'd2 : wc_rawsize;
assign wc_burst = wc_bus[59:58];
// =======================================================================
// Write Response Path Processing
// =======================================================================
// ============================================
// Write Response header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  ws_hdr            = {24{1'b0}};
  // Assign over the various fields
  ws_hdr[3:0]  = wc_qos;                                                        // loopback QoS from write command
  ws_hdr[6:4]  = wc_sid;                                                        // loopback SID from write command to DID
  ws_hdr[7]  = 1'b1;                                                            // SoT: not supporting fragmentation yet
  ws_hdr[8]  = 1'b1;                                                            // EoT: not supporting fragmentation yet
  ws_hdr[14:9]  = 6'd3;                                                         // Read command
  ws_hdr[17:15]  = wc_did;                                                      // loopback DID from wrtie command to SID
  ws_hdr[19:18]   = wc_id;
  ws_hdr[23:20] = pslverrWr_4bit;
end

// declare the state parameters for read
parameter S_RC_HDR = 2'd0;
parameter S_RDS_WAIT = 2'd1;
parameter S_RDS_HDR = 2'd2;
parameter S_RDS_PLD = 2'd3;
// ============================================
// Write Response header pslverr latching
// ============================================
assign setWrError = (int_psel &&  int_penable && int_pwrite && int_pready && int_pslverr);
assign clrWrError = (wr_state == 2'd0);
assign pslverrWr_4bit = (setWrError || pslverrWr_latch) ? 4'd2 : 4'd0;
// Latching valid pslverr
always_ff @(posedge clk, negedge frst_n)
begin
  if (!frst_n)
    pslverrWr_latch <= #1ps 1'd0;
  else if (clrWrError || setWrError)
    pslverrWr_latch <= #1ps pslverrWr_latch_nxt;
end

always_comb
begin
  pslverrWr_latch_nxt = pslverrWr_latch;
  // Reset the latched signal for each data phase
  if (clrWrError)
    pslverrWr_latch_nxt = 1'b0;
  // Set the latched signal if performing data phase and slave error is asserted
  else if (setWrError)
    pslverrWr_latch_nxt = 1'b1;
end

// ============================================
// Read Response header pslverr latching
// ============================================
assign setRdError = (int_psel &&  int_penable && !int_pwrite && int_pready && int_pslverr) && (rd_state == S_RDS_WAIT);
assign clrRdError = (rd_state == 2'd0);
assign pslverrRd_4bit = (setRdError || pslverrRd_latch) ? 4'd2 : 4'd0;
// Latching valid pslverr
always_ff @(posedge clk, negedge frst_n)
begin
  if (!frst_n)
    pslverrRd_latch <= #1ps 1'd0;
  else if (clrRdError || setRdError)
    pslverrRd_latch <= #1ps pslverrRd_latch_nxt;
end

always_comb
begin
  pslverrRd_latch_nxt = pslverrRd_latch;
  // Reset the latched signal for each data phase
  if (clrRdError)
    pslverrRd_latch_nxt = 1'b0;
  // Set the latched signal if performing data phase and slave error is asserted
  else if (setRdError)
    pslverrRd_latch_nxt = 1'b1;
end

// =======================================================================
// Read Processing
// =======================================================================
// Current Read Flit Count
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rc_cnt <= #1ps 1'd0;
  else if (rc_cnt_en)
    rc_cnt <= #1ps rc_cnt_nxt;
end

assign prdata = int_prdata;
assign pslverr_w = int_pslverr;
// Read State Machine State
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rd_state <= #1ps S_RC_HDR;
  else if (rd_state_en)
    rd_state <= #1ps rd_state_nxt;
end

// Read Command Packing Buffer
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rc_buf[0] <= #1ps {60{1'b0}};
    end
  else
    begin
      if (rc_buf_en[0])
        rc_buf[0] <= #1ps if1_flitdata;
    end
end

assign rc_buf_en = rc_buf_we << rc_cnt;
// ============================================
// Read Data + Status flit sequencer
// ============================================
always_comb
begin
  // Defaults
  rd_state_nxt  = rd_state;
  rc_cnt_nxt    = rc_cnt;
  ir0_req       = 1'b0;
  ir0_sop       = 1'b0;
  ir0_eop       = 1'b0;
  ir0_flitdata  = {34{1'b0}};
  rds_transinfo_we = 1'b0;
  if1_ready     = 1'b0;
  rf_ready      = 1'b0;
  // Write enables
  rd_state_en   = 1'b0;
  rc_cnt_en     = 1'b0;
  rc_buf_we     = 1'b0;
  int_arvalid  = 1'b0;
  case (rd_state)
    S_RC_HDR:
      begin
        if1_ready    = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if1_req)
          begin
            // Header transmission is complete
            if (rc_cnt == 1'd0)
              begin
                int_arvalid  = 1'b1;
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rc_buf_we    = 1'b1;
                rds_transinfo_we = 1'b1;
                rd_state_nxt = S_RDS_WAIT;
                rd_state_en   = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                rc_buf_we    = 1'b1;
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
   S_RDS_WAIT:
   begin
    if (int_pready && int_penable && !int_pwrite)
    begin
        rd_state_nxt = S_RDS_HDR;
        rd_state_en  = 1'b1;
    end
   end
   S_RDS_HDR:
      begin
        ir0_req   = 1'd1;
        ir0_sop   = (rc_cnt == 1'd0);
        case(rc_cnt)
          1'd0: ir0_flitdata = rds_hdr[33:0];
          1'd1: ir0_flitdata = rds_hdr[67:34];
          default: ir0_flitdata = {34{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir0_req && ir0_ready)
          begin
            // Complete header is done
            if (rc_cnt == 1'd1)
              begin
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rd_state_nxt = S_RDS_PLD;
                rd_state_en   = 1'b1;
              end
            else
              begin
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
    S_RDS_PLD:
      begin
        ir0_req       = rf_req;
        ir0_eop       = rf_eop;
        ir0_flitdata  = rf_flitdata;
        rf_ready      = ir0_ready;
        if (rf_req && rf_eop && ir0_ready)
          begin
            rd_state_nxt = S_RC_HDR;
            rd_state_en   = 1'b1;
          end
      end
  endcase
end

always_ff @(posedge rcclk) assert ( (frst_n===1'b0) || (int_arvalid == 1'b0) || (rc_burst != 2'b00) || ({{(32-3){1'b0}},rc_plen} <= (32<<1) ) ) else $error("ERROR usb4_tc_noc_apbtea4 : %0t : Read data burst request is larger than TEA can handle. Read data burst size(rplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,rc_plen,(32<<1) );
usb4_tc_noc_apbtea4_rdpack rdpack (
  .clk(rdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .tr_req(rds_transinfo_we),                                                    // i:1
  .tr_rdy(rds_transinfo_rdy),                                                   // o:1
  .tr_size(rc_size),                                                            // i:3
  .tr_burst(rc_burst),                                                          // i:2
  .tr_addrlsb(rc_addr[11:0]),                                                   // i:12
  .tr_plen(rc_plen),                                                            // i:3
  .r_req(rd_req),                                                               // o:1
  .r_last(rd_last),                                                             // o:1
  .r_data(prdata),                                                              // i:32
  .r_slverr(pslverr_w),                                                         // i:1
  .r_ready(rd_ready),                                                           // i:1
  .f_req(rf_req),                                                               // o:1
  .f_eop(rf_eop),                                                               // o:1
  .f_flitdata(rf_flitdata),                                                     // o:34
  .f_ready(rf_ready),                                                           // i:1
  .tr_addrlsb_out(rc_addr_pack)                                                 // o:12
);
// Create incoming rc bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rc_bus[59:0] = (rd_state == S_RC_HDR) ? if1_flitdata : rc_buf[0];
// assign rc.bus = {$rcBusStr};
// Read Command Signal Unpacking
assign rc_sid = rc_bus[17:15];
assign rc_did = rc_bus[6:4];
assign rc_id = rc_bus[19:18];
assign rc_addr = rc_bus[54:23];
assign rc_qos = rc_bus[3:0];
assign rc_plen = rc_bus[22:20];
assign rc_prot = 3'd0;
assign rc_rawsize = rc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign rc_size = Narrow_Req ? ((rc_rawsize < 3'd2) ? rc_rawsize : 3'd2) : ((rc_rawsize > 3'd2) ? 3'd2 : rc_rawsize);
assign rc_burst = rc_bus[59:58];
assign Narrow_Req = rc_rawsize < 3'd2;
// ============================================
// Read Data + Status Header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  rds_hdr            = {68{1'b0}};
  // Assign over the various fields
  rds_hdr[3:0]  = rc_qos;                                                       // loopback QoS from write command
  rds_hdr[6:4]  = rc_sid;                                                       // loopback SID from write command to DID
  rds_hdr[7]  = 1'b1;                                                           // SoT: not supporting fragmentation yet
  rds_hdr[8]  = 1'b1;                                                           // EoT: not supporting fragmentation yet
  rds_hdr[14:9]  = 6'd1;                                                        // Read data / status
  rds_hdr[17:15]  = rc_did;                                                     // loopback DID from wrtie command to SID
  rds_hdr[19:18]   = rc_id;
  rds_hdr[22:20] = rc_plen;
  rds_hdr[30:23]  = (rc_burst==2'd2) ? 8'(rc_addr[11:0] >> rc_size) : rc_addr[7:0];
  rds_hdr[33:31]  = rc_size;
  rds_hdr[35:34] = rc_burst;
end

// Arbitrate between read and write state machines for use of APB interface
parameter S_PSEL = 2'd0;
parameter S_PWEN = 2'd1;
parameter S_PREN = 2'd2;
parameter S_PRDATA = 2'd3;
// APB State Machine State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_state <= #1ps S_PSEL;
  else if (apb_state_en)
    apb_state <= #1ps apb_state_nxt;
end

// Read / Write Arbiter State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_wrarb <= #1ps 1'd0;
  else if (apb_wrarb_en)
    apb_wrarb <= #1ps apb_wrarb_nxt;
end

// For multiple targets and when both rd and wr are active
always_comb
begin
  int_psel      = 1'b0;
  int_pwrite    = 1'b0;
  int_penable   = 1'b0;
  int_paddr     = {18{1'b0}};
  int_pwdata    = {32{1'b0}};
  int_pstrb     = {4{1'b0}};
  int_pprot     = 3'd0;
  apb_state_nxt = apb_state;
  apb_state_en  = 1'b0;
  apb_wrarb_nxt = apb_wrarb;
  apb_wrarb_en  = 1'b0;
  wr_ready      = 1'b0;
  rd_ready      = 1'b0;
  case (apb_state)
    S_PSEL:
      begin
        if (wr_req && (!rd_req || apb_wrarb))
          begin
            int_psel      = 1'b1;
            int_paddr     = {wc_addr[17:12],wc_addr_unpack};
            int_pwrite    = 1'b1;
            int_pwdata    = wr_data;
            int_pstrb     = wr_strb;
            int_pprot     = wc_prot;
            apb_state_nxt = S_PWEN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b0;
            apb_wrarb_en  = 1'b1;
          end
        else if (rd_req)
          begin
            int_psel      = 1'b1;
            int_paddr     = {rc_addr[17:12],rc_addr_pack};
            int_pprot     = rc_prot;
            apb_state_nxt = S_PREN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b1;
            apb_wrarb_en  = 1'b1;
          end
      end
    S_PWEN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
        int_pwrite  = 1'b1;
        int_paddr   = {wc_addr[17:12],wc_addr_unpack};
        int_pwdata  = wr_data;
        int_pstrb   = wr_strb;
        int_pprot   = wc_prot;
        if (int_pready)
          begin
            wr_ready   = 1'b1;
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
          end
      end
    S_PREN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
            int_paddr     = {rc_addr[17:12],rc_addr_pack};
        int_pprot   = rc_prot;
        if (int_pready)
          begin
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
            rd_ready   = 1'b1;
          end
      end
    // S_PRDATA:
    // begin
    // apb.state.nxt = S_PSEL;
    // apb.state.en  = 1'b1;
    // end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_epipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire     [17:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  output logic           src_pslverr,                                           // Slave error
  // dst
  output logic    [17:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata,                                            // Read data
  input  wire            dst_pslverr                                            // Slave error
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea4_epipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
assign src_pslverr = dst_pslverr;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_epipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea4_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea4_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea4_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea4_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_apbcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_wccg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_wdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_f1cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_rdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_wdunpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wtr_req,
  output logic           wtr_rdy,
  input  wire      [2:0] wtr_size,                                              // Transfer size per data phase
  input  wire      [1:0] wtr_burst,                                             // Burst addressing mode
  input  wire     [11:0] wtr_addrlsb,                                           // 12 LSBs of address
  input  wire      [2:0] wtr_plen,                                              // Packet length in bytes
  output logic           w_valid,
  output logic    [31:0] w_data,
  output logic     [3:0] w_strb,
  output logic           w_last,
  input  wire            w_ready,
  input  wire            f_req,
  input  wire            f_eop,
  input  wire     [35:0] f_flitdata,
  output logic           f_ready,
  output logic    [11:0] wtr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [2:0] sizeCnvDiv;
logic     [4:0] firstCnt2Wrap;
logic     [7:0] wtr_mask;
logic     [7:0] wtr_mis;
logic    [10:0] firstXferCnt;
logic    [10:0] xferCnt;
logic    [10:0] xferCnt_nxt;
logic     [0:0] xferCnt_en;
logic    [10:0] useXferCnt;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic    [31:0] muxed_w_data;
logic     [3:0] muxed_w_strb;
logic           flitDone;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic     [0:0] haveFlit;
logic     [0:0] haveFlit_nxt;
logic     [0:0] haveFlit_en;
logic    [35:0] flitData;
logic    [35:0] flitData_nxt;
logic     [0:0] flitData_en;
logic           flitValid;
logic    [11:0] lower_baddr;
logic    [11:0] upper_baddr;
logic    [11:0] lower_addr;
logic    [11:0] upper_addr;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
logic    [11:0] saddr;
logic     [2:0] splen;
// Extracted from packet header
// APB W Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},wtr_plen} - 1'b1;                                    // We only care about 8 bits of address for our word indexing
assign wrapToAddr = wtr_addrlsb[7:0] & ~bamask;                                 // This is the address offset we wrap to
assign wrapIndex = wtr_addrlsb >> wtr_size;
assign sizeCnvDiv = wtr_plen >> wtr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign wtr_mask = (8'b1<<wtr_size) - 1'b1;
assign wtr_mis = wtr_addrlsb[7:0] & wtr_mask;
assign firstXferCnt = (wtr_burst!=2'd1) ? 11'(wtr_plen>>wtr_size) : 11'((16'(wtr_plen)+wtr_mask+wtr_mis)>>wtr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    xferCnt <= #1ps 11'd0;
  else if (xferCnt_en)
    xferCnt <= #1ps xferCnt_nxt;
end

assign useXferCnt = xferCnt;
always_comb
begin
  xferCnt_nxt = xferCnt;
  xferCnt_en  = 1'b0;
  if( newCmd )
    begin
      xferCnt_nxt = firstXferCnt;
      xferCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      xferCnt_nxt = useXferCnt - 1'd1;
      xferCnt_en  = 1'b1;
    end
end

assign wtr_rdy = ~trInPkt;
assign newCmd = wtr_req && wtr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = w_valid && w_ready;
assign f_ready = ~haveFlit || flitDone;
assign w_valid = flitValid;
assign w_last = w_valid && useXferCnt==11'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps wtr_burst;
end

assign use_tr_burst = held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps wtr_size;
end

assign use_tr_size = held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( busWriteValid && w_last )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> wtr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (wtr_addrlsb[7:0] & 8'd3) >> wtr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( w_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone;
assign muxed_w_data[7:0] = flitData[7:0];
assign muxed_w_strb[3:0] = flitData[35:32];
assign muxed_w_data[15:8] = flitData[15:8];
assign muxed_w_data[23:16] = flitData[23:16];
assign muxed_w_data[31:24] = flitData[31:24];
assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    haveFlit <= #1ps 1'd0;
  else if (haveFlit_en)
    haveFlit <= #1ps haveFlit_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitData <= #1ps {36{1'b0}};
  else if (flitData_en)
    flitData <= #1ps flitData_nxt;
end

assign flitValid = haveFlit;
always_comb
begin
  haveFlit_nxt   = haveFlit;
  haveFlit_en    = 1'b0;
  flitData_nxt   = flitData;
  flitData_en    = 1'b0;
  if( flitWriteValid )
    begin
      haveFlit_nxt   = 1'b1;
      haveFlit_en    = 1'b1;
      flitData_en    = 1'b1;
      flitData_nxt   = f_flitdata;
    end
  else if( flitDone )
    begin
      haveFlit_nxt   = 1'b0;
      haveFlit_en    = 1'b1;
    end
end

assign w_data[7:0] = (w_valid && wrMask[0]) ? muxed_w_data[7:0] : 8'd0;
assign w_data[15:8] = (w_valid && wrMask[1]) ? muxed_w_data[15:8] : 8'd0;
assign w_data[23:16] = (w_valid && wrMask[2]) ? muxed_w_data[23:16] : 8'd0;
assign w_data[31:24] = (w_valid && wrMask[3]) ? muxed_w_data[31:24] : 8'd0;
assign w_strb = w_valid ? muxed_w_strb & wrMask : 4'd0;
assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  addrlsb_nxt   = addrlsb;
  // Write enables
  addrlsb_en    = 1'b0;
  if (newCmd)
    begin
      addrlsb_nxt = wtr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred from packing FIFO
  else if (busWriteValid)
    begin
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps wtr_addrlsb;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps wtr_plen;
end

assign wtr_addrlsb_out = !(newCmd) ? addrlsb : wtr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea4_rdpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            tr_req,
  output logic           tr_rdy,
  input  wire      [2:0] tr_size,
  input  wire      [1:0] tr_burst,
  input  wire     [11:0] tr_addrlsb,
  input  wire      [2:0] tr_plen,
  output logic           r_req,
  output logic           r_last,
  input  wire     [31:0] r_data,
  input  wire            r_slverr,
  input  wire            r_ready,
  output logic           f_req,
  output logic           f_eop,
  output logic    [33:0] f_flitdata,
  input  wire            f_ready,
  output logic    [11:0] tr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [4:0] firstCnt2Wrap;
logic     [2:0] sizeCnvDiv;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [0:0] heldFlitDone;
logic     [0:0] heldEop;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isNarrow;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic           flitDone;
logic           useBusWdCnt;
logic    [33:0] flitWd;
logic    [33:0] flitWd_nxt;
logic     [0:0] flitWd_en;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] lower_baddr;                                                    // Lower burst address
logic    [11:0] upper_baddr;                                                    // Upper burst address
logic    [11:0] lower_addr;                                                     // Lower element address
logic    [11:0] upper_addr;                                                     // Upper element address
logic    [11:0] esize_minus_first_offset;
logic    [11:0] first_offset;
logic     [2:0] raw_wcnt;
logic     [2:0] wcnt;
logic    [11:0] saddr;
logic     [2:0] wplen;
logic     [2:0] wplen_nxt;
logic     [0:0] wplen_en;
logic     [2:0] splen;
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
// Extracted from AXI AW Channel
// APB R Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},tr_plen} - 1'b1;                                     // We only care about 8 bits of address for our word indexing
assign wrapToAddr = tr_addrlsb[7:0] & ~bamask;                                  // This is the address offset we wrap to
assign wrapIndex = tr_addrlsb >> tr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign sizeCnvDiv = tr_plen >> tr_size;
assign tr_rdy = ~trInPkt;
assign f_flitdata = flitWd;
assign f_req = heldFlitDone;
assign f_eop = heldEop;
assign r_req = trInPkt_nxt && (!heldFlitDone || flitWriteValid);
assign newCmd = tr_req && tr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = r_ready && r_req;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldFlitDone <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldFlitDone <= #1ps flitDone;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldEop <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldEop <= #1ps flitDone && r_last;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps tr_burst;
end

assign use_tr_burst = (newCmd) ? tr_burst : held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps tr_size;
end

assign use_tr_size = (newCmd) ? tr_size : held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isNarrow = use_tr_size<3'd2;
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( flitWriteValid && f_eop )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> tr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = (newCmd) ? subBusWdCntWrap_nxt : subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = newCmd ? firstCnt2Wrap : cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (tr_addrlsb[7:0] & 8'd3) >> tr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = (newCmd) ? firstSubBusWdCnt[1:0] : subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( r_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone || (isNarrow && busWriteValid);
assign useBusWdCnt = 1'b0;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitWd <= #1ps {34{1'b0}};
  else if (flitWd_en)
    flitWd <= #1ps flitWd_nxt;
end

assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_comb
begin
  // First, assign the bus word to every possible flit word slot
  flitWd_nxt = flitWriteValid ? {34{1'b0}} : flitWd;
  // Start out with nothing enabled
  flitWd_en = flitWriteValid ? 1'b1 : 1'b0;
  // Now enable any bytes that are being written this cycle
  if( busWriteValid )
    begin
      if( useBusWdCnt == 1'd0 )
        begin
          if( wrMask[0] )
            begin
              flitWd_nxt[7:0] = r_data[7:0];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[1] )
            begin
              flitWd_nxt[15:8] = r_data[15:8];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[2] )
            begin
              flitWd_nxt[23:16] = r_data[23:16];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[3] )
            begin
              flitWd_nxt[31:24] = r_data[31:24];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
        end
    end
end

assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
assign esize_minus_first_offset = esize - first_offset;
assign first_offset = addrlsb & amask;
assign raw_wcnt = (held_tr_burst == 2'd1) ? esize_minus_first_offset[2:0] : esize[2:0];
assign wcnt = (raw_wcnt > wplen) ? wplen : raw_wcnt;
assign r_last = (wcnt >= wplen);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps tr_addrlsb;
end

// Write remaining packet length and address LSB tracking flops
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    wplen <= #1ps 3'd0;
  else if (wplen_en)
    wplen <= #1ps wplen_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps tr_plen;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  wplen_nxt   = wplen;
  addrlsb_nxt = addrlsb;
  wplen_en    = 1'b0;
  addrlsb_en  = 1'b0;
  if (tr_req && tr_rdy)
    begin
      wplen_nxt   = tr_plen;
      wplen_en    = 1'b1;
      addrlsb_nxt = tr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred to packing FIFO
  else if (busWriteValid)
    begin
      wplen_en    = 1'b1;
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            wplen_nxt   = wplen - wcnt;
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            wplen_nxt   = wplen   - wcnt;
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            wplen_nxt   = wplen      - wcnt;
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            wplen_nxt   = wplen;
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

assign tr_addrlsb_out = !(newCmd) ? addrlsb : tr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5 (
  input  wire            clk,
  input  wire            rst_n,
  // t
  output logic     [9:0] t_paddr,                                               // Address
  output logic           t_psel,                                                // Select
  output logic           t_penable,                                             // Enable
  output logic           t_pwrite,                                              // Write not read
  output logic    [31:0] t_pwdata,                                              // Write data
  output logic     [3:0] t_pstrb,                                               // Write strobes
  input  wire            t_pready,                                              // Ready
  input  wire     [31:0] t_prdata,                                              // Read data
  // f0
  input  wire            f0_activity,                                           // Upcoming activity indicator
  input  wire            f0_req,                                                // Flit transfer request
  input  wire            f0_sop,                                                // Start of packet indicator
  input  wire            f0_eop,                                                // End of packet indicator
  input  wire     [35:0] f0_flitdata,                                           // Flit data
  output logic           f0_ready,                                              // Flit transfer ready
  // f1
  input  wire            f1_activity,                                           // Upcoming activity indicator
  input  wire            f1_req,                                                // Flit transfer request
  input  wire            f1_sop,                                                // Start of packet indicator
  input  wire            f1_eop,                                                // End of packet indicator
  input  wire     [59:0] f1_flitdata,                                           // Flit data
  output logic           f1_ready,                                              // Flit transfer ready
  // r0
  output logic           r0_activity,                                           // Upcoming activity indicator
  output logic           r0_req,                                                // Flit transfer request
  output logic           r0_sop,                                                // Start of packet indicator
  output logic           r0_eop,                                                // End of packet indicator
  output logic    [33:0] r0_flitdata,                                           // Flit data
  input  wire            r0_ready,                                              // Flit transfer ready
  // r1
  output logic           r1_activity,                                           // Upcoming activity indicator
  output logic           r1_req,                                                // Flit transfer request
  output logic           r1_sop,                                                // Start of packet indicator
  output logic           r1_eop,                                                // End of packet indicator
  output logic    [23:0] r1_flitdata,                                           // Flit data
  input  wire            r1_ready                                               // Flit transfer ready
);

logic     [9:0] int_paddr;                                                      // Address
logic           int_psel;                                                       // Select
logic           int_penable;                                                    // Enable
logic           int_pwrite;                                                     // Write not read
logic    [31:0] int_pwdata;                                                     // Write data
logic     [3:0] int_pstrb;                                                      // Write strobes
logic           int_pready;                                                     // Ready
logic    [31:0] int_prdata;                                                     // Read data
logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic           wr_req;
logic           wr_ready;
logic           wr_last;
logic    [31:0] wr_data;
logic     [3:0] wr_strb;
logic           wc_buf_we;
logic    [71:0] wc_bus;
logic     [2:0] wc_sid;
logic     [2:0] wc_did;
logic     [1:0] wc_id;
logic    [31:0] wc_addr;
logic     [7:0] wc_len;
logic     [2:0] wc_rawsize;
logic     [2:0] wc_size;
logic     [1:0] wc_burst;
logic     [3:0] wc_qos;
logic     [2:0] wc_plen;
logic     [2:0] wc_prot;
logic           wcd_transinfo_en;
logic           wcd_transinfo_rdy;
logic           wf_req;
logic           wf_eop;
logic    [35:0] wf_flitdata;
logic           wf_ready;
logic    [23:0] ws_hdr;
logic           int_awvalid;
logic    [67:0] rds_hdr;
logic           rd_req;
logic           rd_ready;
logic           rd_last;
logic           rc_buf_we;
logic    [59:0] rc_bus;
logic     [2:0] rc_sid;
logic     [2:0] rc_did;
logic     [1:0] rc_id;
logic    [31:0] rc_addr;
logic     [2:0] rc_rawsize;
logic     [2:0] rc_size;
logic     [1:0] rc_burst;
logic     [3:0] rc_qos;
logic     [2:0] rc_plen;
logic     [2:0] rc_prot;
logic           rf_req;
logic           rf_eop;
logic    [33:0] rf_flitdata;
logic           rf_ready;
logic           rds_transinfo_we;
logic           rds_transinfo_rdy;
logic           int_arvalid;
logic    [11:0] wc_addr_unpack;
logic    [11:0] rc_addr_pack;
logic     [2:0] int_pprot;
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           apbclk;
logic           apbclkAct;
logic           int_apbactivity;
logic           wcclk;
logic           wcclkAct;
wire            int_awactivity;
logic           wdclk;
logic           wdclkAct;
logic           int_wactivity;
logic           rcclk;
logic           rcclkAct;
logic           int_aractivity;
logic           rdclk;
logic           rdclkAct;
logic           rdclkEn;
logic           wrDone;
logic     [0:0] wr_cnt;
logic     [0:0] wr_cnt_nxt;
logic     [0:0] wr_cnt_en;
logic     [1:0] wr_state;
logic     [1:0] wr_state_nxt;
logic     [0:0] wr_state_en;
logic    [35:0] wc_buf [1:0];
logic     [1:0] wc_buf_en;
logic           int_pslverr;
logic     [0:0] rc_cnt;
logic     [0:0] rc_cnt_nxt;
logic     [0:0] rc_cnt_en;
logic           pslverr_w;
logic    [31:0] prdata;
logic     [1:0] rd_state;
logic     [1:0] rd_state_nxt;
logic     [0:0] rd_state_en;
logic    [59:0] rc_buf [0:0];
logic     [0:0] rc_buf_en;
logic           Narrow_Req;
logic     [1:0] apb_state;
logic     [1:0] apb_state_nxt;
logic     [0:0] apb_state_en;
logic     [0:0] apb_wrarb;
logic     [0:0] apb_wrarb_nxt;
logic     [0:0] apb_wrarb_en;
// ========================================================================//
// Parameter Declarations
// ========================================================================//
// ========================================================================//
// Process parameters and create local derived variables
// ========================================================================//
// ========================================================================//
// Define module I/O
// ========================================================================//
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// APB Target Interface(s) (APB manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// Egress APB Pipeline Component
usb4_tc_noc_apbtea5_epipe epipe (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .src_paddr(int_paddr),                                                        // i:10
  .src_psel(int_psel),                                                          // i:1
  .src_penable(int_penable),                                                    // i:1
  .src_pwrite(int_pwrite),                                                      // i:1
  .src_pwdata(int_pwdata),                                                      // i:32
  .src_pstrb(int_pstrb),                                                        // i:4
  .src_pready(int_pready),                                                      // o:1
  .src_prdata(int_prdata),                                                      // o:32
  .dst_paddr(t_paddr),                                                          // o:10
  .dst_psel(t_psel),                                                            // o:1
  .dst_penable(t_penable),                                                      // o:1
  .dst_pwrite(t_pwrite),                                                        // o:1
  .dst_pwdata(t_pwdata),                                                        // o:32
  .dst_pstrb(t_pstrb),                                                          // o:4
  .dst_pready(t_pready),                                                        // i:1
  .dst_prdata(t_prdata)                                                         // i:32
);
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea5_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f0_activity),                                                   // i:1
  .src_req(f0_req),                                                             // i:1
  .src_sop(f0_sop),                                                             // i:1
  .src_eop(f0_eop),                                                             // i:1
  .src_flitdata(f0_flitdata),                                                   // i:36
  .src_ready(f0_ready),                                                         // o:1
  .dst_activity(if0_activity),                                                  // o:1
  .dst_req(if0_req),                                                            // o:1
  .dst_sop(if0_sop),                                                            // o:1
  .dst_eop(if0_eop),                                                            // o:1
  .dst_flitdata(if0_flitdata),                                                  // o:36
  .dst_ready(if0_ready)                                                         // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_apbtea5_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f1_activity),                                                   // i:1
  .src_req(f1_req),                                                             // i:1
  .src_sop(f1_sop),                                                             // i:1
  .src_eop(f1_eop),                                                             // i:1
  .src_flitdata(f1_flitdata),                                                   // i:60
  .src_ready(f1_ready),                                                         // o:1
  .dst_activity(if1_activity),                                                  // o:1
  .dst_req(if1_req),                                                            // o:1
  .dst_sop(if1_sop),                                                            // o:1
  .dst_eop(if1_eop),                                                            // o:1
  .dst_flitdata(if1_flitdata),                                                  // o:60
  .dst_ready(if1_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea5_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir0_activity),                                                  // i:1
  .src_req(ir0_req),                                                            // i:1
  .src_sop(ir0_sop),                                                            // i:1
  .src_eop(ir0_eop),                                                            // i:1
  .src_flitdata(ir0_flitdata),                                                  // i:34
  .src_ready(ir0_ready),                                                        // o:1
  .dst_activity(r0_activity),                                                   // o:1
  .dst_req(r0_req),                                                             // o:1
  .dst_sop(r0_sop),                                                             // o:1
  .dst_eop(r0_eop),                                                             // o:1
  .dst_flitdata(r0_flitdata),                                                   // o:34
  .dst_ready(r0_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_apbtea5_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir1_activity),                                                  // i:1
  .src_req(ir1_req),                                                            // i:1
  .src_sop(ir1_sop),                                                            // i:1
  .src_eop(ir1_eop),                                                            // i:1
  .src_flitdata(ir1_flitdata),                                                  // i:24
  .src_ready(ir1_ready),                                                        // o:1
  .dst_activity(r1_activity),                                                   // o:1
  .dst_req(r1_req),                                                             // o:1
  .dst_sop(r1_sop),                                                             // o:1
  .dst_eop(r1_eop),                                                             // o:1
  .dst_flitdata(r1_flitdata),                                                   // o:24
  .dst_ready(r1_ready)                                                          // i:1
);
// =======================================================================
// Signal declarations
// =======================================================================
// Write Command + Data Sequencer Signals
// Write Command Signals
// Write Response Fields
// Read Data + Status fields
// Read Data + Status Flit Sequencer Signals
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea5_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign int_apbactivity = int_awactivity || int_aractivity;
usb4_tc_noc_apbtea5_apbcg apbcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_apbactivity),                                                      // i:1
  .clkOut(apbclk),                                                              // o:1
  .isActive(apbclkAct)                                                          // o:1
);
assign int_awactivity = if0_activity || if0_req || int_awvalid || ir1_req || wr_req;
usb4_tc_noc_apbtea5_wccg wccg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_awactivity),                                                       // i:1
  .clkOut(wcclk),                                                               // o:1
  .isActive(wcclkAct)                                                           // o:1
);
assign int_wactivity = if0_activity || if0_req || !wcd_transinfo_rdy || int_awvalid;
usb4_tc_noc_apbtea5_wdcg wdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_wactivity),                                                        // i:1
  .clkOut(wdclk),                                                               // o:1
  .isActive(wdclkAct)                                                           // o:1
);
assign ir1_activity = ir1_req;
assign int_aractivity = if1_activity || if1_req || ir0_req || rd_req;
usb4_tc_noc_apbtea5_f1cg f1cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(int_aractivity),                                                       // i:1
  .clkOut(rcclk),                                                               // o:1
  .isActive(rcclkAct)                                                           // o:1
);
assign ir0_activity = ir0_req;
assign rdclkEn = ir0_activity || if1_activity || if1_req || !rds_transinfo_rdy;
usb4_tc_noc_apbtea5_rdcg rdcg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(rdclkEn),                                                              // i:1
  .clkOut(rdclk),                                                               // o:1
  .isActive(rdclkAct)                                                           // o:1
);
// =======================================================================
// Write Processing
// =======================================================================
assign wrDone = wr_last && int_penable && int_pwrite && int_pready;
parameter S_WR_HDR = 2'd0;
parameter S_WR_DATA = 2'd1;
parameter S_WR_WAIT = 2'd2;
parameter S_WR_STS = 2'd3;
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign wc_bus[35:0] = wc_buf[0];
assign wc_bus[71:36] = ((wr_state == 2'b00) && (wr_cnt >= 1'd1)) ? if0_flitdata : wc_buf[1];
// Current Flit Count
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_cnt <= #1ps 1'd0;
  else if (wr_cnt_en)
    wr_cnt <= #1ps wr_cnt_nxt;
end

// Write State Machine State
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    wr_state <= #1ps S_WR_HDR;
  else if (wr_state_en)
    wr_state <= #1ps wr_state_nxt;
end

// Write Command Packing Buffer
always_ff @(posedge wcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      wc_buf[0] <= #1ps {36{1'b0}};
      wc_buf[1] <= #1ps {36{1'b0}};
    end
  else
    begin
      if (wc_buf_en[0])
        wc_buf[0] <= #1ps if0_flitdata;
      if (wc_buf_en[1])
        wc_buf[1] <= #1ps if0_flitdata;
    end
end

assign wc_buf_en = wc_buf_we << wr_cnt;
always_comb
begin
  // Defaults
  if0_ready    = 1'b0;
  ir1_req      = 1'b0;
  ir1_sop      = 1'b0;
  ir1_eop      = 1'b0;
  ir1_flitdata = {24{1'b0}};
  wr_cnt_nxt   = wr_cnt;
  wr_state_nxt = wr_state;
  wcd_transinfo_en = 1'b0;
  wf_req       = 1'b0;
  wf_eop       = 1'b0;
  wf_flitdata  = {36{1'b0}};
  // Write enables
  wc_buf_we    = 1'b0;
  wr_cnt_en    = 1'b0;
  wr_state_en  = 1'b0;
  int_awvalid   = 1'b0;
  case (wr_state)
    S_WR_HDR:
      begin
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_req)
          begin
            if0_ready    = 1'b1;
            // Header transmission is complete
            if (wr_cnt == 1'd1)
              begin
                int_awvalid = wcd_transinfo_rdy;
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wc_buf_we    = 1'b1;
                wcd_transinfo_en = 1'b1;
                wr_state_nxt = S_WR_DATA;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
                wc_buf_we  = 1'b1;
              end
          end
      end
   S_WR_DATA:
      begin
        wf_req      = if0_req;
        wf_eop      = if0_eop;
        wf_flitdata = if0_flitdata;
        if0_ready   = wf_ready;
        if (if0_req && wf_ready && if0_eop)
          begin
            wr_state_nxt = S_WR_WAIT;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_WAIT:
      begin
        if (wr_req && wr_ready && wr_last)
          begin
            wr_state_nxt = S_WR_STS;
            wr_state_en  = 1'b1;
          end
      end
    S_WR_STS:
      begin
        ir1_req   = 1'b1;
        ir1_sop   = (wr_cnt == 1'd0);
        ir1_eop   = (wr_cnt == 1'd0);
        case(wr_cnt)
          1'd0: ir1_flitdata = ws_hdr[23:0];
          default: ir1_flitdata = {24{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_ready)
          begin
            // Header transmission is complete
            if (wr_cnt == 1'd0)
              begin
                wr_cnt_nxt   = 1'd0;
                wr_cnt_en    = 1'b1;
                wr_state_nxt = S_WR_HDR;
                wr_state_en  = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                wr_cnt_nxt = wr_cnt + 1'd1;
                wr_cnt_en  = 1'b1;
              end
          end
      end
  endcase
end

 always_ff @(posedge wcclk) assert ( (frst_n===1'b0) || (int_awvalid == 1'b0) || (wc_burst != 2'b00) || ( {{(32-3){1'b0}},wc_plen} <= (32<<1) )) else $error("ERROR usb4_tc_noc_apbtea5 : %0t : Write data burst request is larger than TEA can handle. Write data burst size(wplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,wc_plen,(32<<1) );
usb4_tc_noc_apbtea5_wdunpack wdunpack (
  .clk(wdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .wtr_req(wcd_transinfo_en),                                                   // i:1
  .wtr_rdy(wcd_transinfo_rdy),                                                  // o:1
  .wtr_size(wc_size),                                                           // i:3
  .wtr_burst(wc_burst),                                                         // i:2
  .wtr_addrlsb(wc_addr[11:0]),                                                  // i:12
  .wtr_plen(wc_plen),                                                           // i:3
  .w_valid(wr_req),                                                             // o:1
  .w_data(wr_data),                                                             // o:32
  .w_strb(wr_strb),                                                             // o:4
  .w_last(wr_last),                                                             // o:1
  .w_ready(wr_ready),                                                           // i:1
  .f_req(wf_req),                                                               // i:1
  .f_eop(wf_eop),                                                               // i:1
  .f_flitdata(wf_flitdata),                                                     // i:36
  .f_ready(wf_ready),                                                           // o:1
  .wtr_addrlsb_out(wc_addr_unpack)                                              // o:12
);
// Write Command + Data Signal Unpacking
assign wc_sid = wc_bus[17:15];
assign wc_did = wc_bus[6:4];
assign wc_id = wc_bus[19:18];
assign wc_addr = wc_bus[54:23];
assign wc_qos = wc_bus[3:0];
assign wc_plen = wc_bus[22:20];
assign wc_prot = 3'd0;
assign wc_rawsize = wc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign wc_size = (wc_rawsize > 3'd2) ? 3'd2 : wc_rawsize;
assign wc_burst = wc_bus[59:58];
// =======================================================================
// Write Response Path Processing
// =======================================================================
// ============================================
// Write Response header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  ws_hdr            = {24{1'b0}};
  // Assign over the various fields
  ws_hdr[3:0]  = wc_qos;                                                        // loopback QoS from write command
  ws_hdr[6:4]  = wc_sid;                                                        // loopback SID from write command to DID
  ws_hdr[7]  = 1'b1;                                                            // SoT: not supporting fragmentation yet
  ws_hdr[8]  = 1'b1;                                                            // EoT: not supporting fragmentation yet
  ws_hdr[14:9]  = 6'd3;                                                         // Read command
  ws_hdr[17:15]  = wc_did;                                                      // loopback DID from wrtie command to SID
  ws_hdr[19:18]   = wc_id;
end

// declare the state parameters for read
parameter S_RC_HDR = 2'd0;
parameter S_RDS_WAIT = 2'd1;
parameter S_RDS_HDR = 2'd2;
parameter S_RDS_PLD = 2'd3;
assign int_pslverr = 1'd0;
// =======================================================================
// Read Processing
// =======================================================================
// Current Read Flit Count
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rc_cnt <= #1ps 1'd0;
  else if (rc_cnt_en)
    rc_cnt <= #1ps rc_cnt_nxt;
end

assign prdata = int_prdata;
assign pslverr_w = int_pslverr;
// Read State Machine State
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    rd_state <= #1ps S_RC_HDR;
  else if (rd_state_en)
    rd_state <= #1ps rd_state_nxt;
end

// Read Command Packing Buffer
always_ff @(posedge rcclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rc_buf[0] <= #1ps {60{1'b0}};
    end
  else
    begin
      if (rc_buf_en[0])
        rc_buf[0] <= #1ps if1_flitdata;
    end
end

assign rc_buf_en = rc_buf_we << rc_cnt;
// ============================================
// Read Data + Status flit sequencer
// ============================================
always_comb
begin
  // Defaults
  rd_state_nxt  = rd_state;
  rc_cnt_nxt    = rc_cnt;
  ir0_req       = 1'b0;
  ir0_sop       = 1'b0;
  ir0_eop       = 1'b0;
  ir0_flitdata  = {34{1'b0}};
  rds_transinfo_we = 1'b0;
  if1_ready     = 1'b0;
  rf_ready      = 1'b0;
  // Write enables
  rd_state_en   = 1'b0;
  rc_cnt_en     = 1'b0;
  rc_buf_we     = 1'b0;
  int_arvalid  = 1'b0;
  case (rd_state)
    S_RC_HDR:
      begin
        if1_ready    = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if1_req)
          begin
            // Header transmission is complete
            if (rc_cnt == 1'd0)
              begin
                int_arvalid  = 1'b1;
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rc_buf_we    = 1'b1;
                rds_transinfo_we = 1'b1;
                rd_state_nxt = S_RDS_WAIT;
                rd_state_en   = 1'b1;
              end
            // Continuing header transmission
            else
              begin
                rc_buf_we    = 1'b1;
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
   S_RDS_WAIT:
   begin
    if (int_pready && int_penable && !int_pwrite)
    begin
        rd_state_nxt = S_RDS_HDR;
        rd_state_en  = 1'b1;
    end
   end
   S_RDS_HDR:
      begin
        ir0_req   = 1'd1;
        ir0_sop   = (rc_cnt == 1'd0);
        case(rc_cnt)
          1'd0: ir0_flitdata = rds_hdr[33:0];
          1'd1: ir0_flitdata = rds_hdr[67:34];
          default: ir0_flitdata = {34{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir0_req && ir0_ready)
          begin
            // Complete header is done
            if (rc_cnt == 1'd1)
              begin
                rc_cnt_nxt   = 1'd0;
                rc_cnt_en    = 1'b1;
                rd_state_nxt = S_RDS_PLD;
                rd_state_en   = 1'b1;
              end
            else
              begin
                rc_cnt_nxt   = rc_cnt + 1'd1;
                rc_cnt_en    = 1'b1;
              end
          end
      end
    S_RDS_PLD:
      begin
        ir0_req       = rf_req;
        ir0_eop       = rf_eop;
        ir0_flitdata  = rf_flitdata;
        rf_ready      = ir0_ready;
        if (rf_req && rf_eop && ir0_ready)
          begin
            rd_state_nxt = S_RC_HDR;
            rd_state_en   = 1'b1;
          end
      end
  endcase
end

always_ff @(posedge rcclk) assert ( (frst_n===1'b0) || (int_arvalid == 1'b0) || (rc_burst != 2'b00) || ({{(32-3){1'b0}},rc_plen} <= (32<<1) ) ) else $error("ERROR usb4_tc_noc_apbtea5 : %0t : Read data burst request is larger than TEA can handle. Read data burst size(rplen)=%d APB TEA data handling capacity=%d Burst=FIXED",$time,rc_plen,(32<<1) );
usb4_tc_noc_apbtea5_rdpack rdpack (
  .clk(rdclk),                                                                  // i:1
  .rst_n(frst_n),                                                               // i:1
  .tr_req(rds_transinfo_we),                                                    // i:1
  .tr_rdy(rds_transinfo_rdy),                                                   // o:1
  .tr_size(rc_size),                                                            // i:3
  .tr_burst(rc_burst),                                                          // i:2
  .tr_addrlsb(rc_addr[11:0]),                                                   // i:12
  .tr_plen(rc_plen),                                                            // i:3
  .r_req(rd_req),                                                               // o:1
  .r_last(rd_last),                                                             // o:1
  .r_data(prdata),                                                              // i:32
  .r_slverr(pslverr_w),                                                         // i:1
  .r_ready(rd_ready),                                                           // i:1
  .f_req(rf_req),                                                               // o:1
  .f_eop(rf_eop),                                                               // o:1
  .f_flitdata(rf_flitdata),                                                     // o:34
  .f_ready(rf_ready),                                                           // i:1
  .tr_addrlsb_out(rc_addr_pack)                                                 // o:12
);
// Create incoming rc bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rc_bus[59:0] = (rd_state == S_RC_HDR) ? if1_flitdata : rc_buf[0];
// assign rc.bus = {$rcBusStr};
// Read Command Signal Unpacking
assign rc_sid = rc_bus[17:15];
assign rc_did = rc_bus[6:4];
assign rc_id = rc_bus[19:18];
assign rc_addr = rc_bus[54:23];
assign rc_qos = rc_bus[3:0];
assign rc_plen = rc_bus[22:20];
assign rc_prot = 3'd0;
assign rc_rawsize = rc_bus[57:55];
// Restrict the size to be less than or equal to the bus width
assign rc_size = Narrow_Req ? ((rc_rawsize < 3'd2) ? rc_rawsize : 3'd2) : ((rc_rawsize > 3'd2) ? 3'd2 : rc_rawsize);
assign rc_burst = rc_bus[59:58];
assign Narrow_Req = rc_rawsize < 3'd2;
// ============================================
// Read Data + Status Header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  rds_hdr            = {68{1'b0}};
  // Assign over the various fields
  rds_hdr[3:0]  = rc_qos;                                                       // loopback QoS from write command
  rds_hdr[6:4]  = rc_sid;                                                       // loopback SID from write command to DID
  rds_hdr[7]  = 1'b1;                                                           // SoT: not supporting fragmentation yet
  rds_hdr[8]  = 1'b1;                                                           // EoT: not supporting fragmentation yet
  rds_hdr[14:9]  = 6'd1;                                                        // Read data / status
  rds_hdr[17:15]  = rc_did;                                                     // loopback DID from wrtie command to SID
  rds_hdr[19:18]   = rc_id;
  rds_hdr[22:20] = rc_plen;
  rds_hdr[30:23]  = (rc_burst==2'd2) ? 8'(rc_addr[11:0] >> rc_size) : rc_addr[7:0];
  rds_hdr[33:31]  = rc_size;
  rds_hdr[35:34] = rc_burst;
end

// Arbitrate between read and write state machines for use of APB interface
parameter S_PSEL = 2'd0;
parameter S_PWEN = 2'd1;
parameter S_PREN = 2'd2;
parameter S_PRDATA = 2'd3;
// APB State Machine State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_state <= #1ps S_PSEL;
  else if (apb_state_en)
    apb_state <= #1ps apb_state_nxt;
end

// Read / Write Arbiter State
always_ff @(posedge apbclk, negedge frst_n)
begin
  if (!frst_n)
    apb_wrarb <= #1ps 1'd0;
  else if (apb_wrarb_en)
    apb_wrarb <= #1ps apb_wrarb_nxt;
end

// For multiple targets and when both rd and wr are active
always_comb
begin
  int_psel      = 1'b0;
  int_pwrite    = 1'b0;
  int_penable   = 1'b0;
  int_paddr     = {10{1'b0}};
  int_pwdata    = {32{1'b0}};
  int_pstrb     = {4{1'b0}};
  int_pprot     = 3'd0;
  apb_state_nxt = apb_state;
  apb_state_en  = 1'b0;
  apb_wrarb_nxt = apb_wrarb;
  apb_wrarb_en  = 1'b0;
  wr_ready      = 1'b0;
  rd_ready      = 1'b0;
  case (apb_state)
    S_PSEL:
      begin
        if (wr_req && (!rd_req || apb_wrarb))
          begin
            int_psel      = 1'b1;
            int_paddr     = wc_addr_unpack[9:0];
            int_pwrite    = 1'b1;
            int_pwdata    = wr_data;
            int_pstrb     = wr_strb;
            int_pprot     = wc_prot;
            apb_state_nxt = S_PWEN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b0;
            apb_wrarb_en  = 1'b1;
          end
        else if (rd_req)
          begin
            int_psel      = 1'b1;
            int_paddr     = rc_addr_pack[9:0];
            int_pprot     = rc_prot;
            apb_state_nxt = S_PREN;
            apb_state_en  = 1'b1;
            apb_wrarb_nxt = 1'b1;
            apb_wrarb_en  = 1'b1;
          end
      end
    S_PWEN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
        int_pwrite  = 1'b1;
        int_paddr   = wc_addr_unpack[9:0];
        int_pwdata  = wr_data;
        int_pstrb   = wr_strb;
        int_pprot   = wc_prot;
        if (int_pready)
          begin
            wr_ready   = 1'b1;
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
          end
      end
    S_PREN:
      begin
        int_psel    = 1'b1;
        int_penable = 1'b1;
            int_paddr     = rc_addr_pack[9:0];
        int_pprot   = rc_prot;
        if (int_pready)
          begin
            apb_state_nxt = S_PSEL;
            apb_state_en  = 1'b1;
            rd_ready   = 1'b1;
          end
      end
    // S_PRDATA:
    // begin
    // apb.state.nxt = S_PSEL;
    // apb.state.en  = 1'b1;
    // end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_epipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire      [9:0] src_paddr,                                             // Address
  input  wire            src_psel,                                              // Select
  input  wire            src_penable,                                           // Enable
  input  wire            src_pwrite,                                            // Write not read
  input  wire     [31:0] src_pwdata,                                            // Write data
  input  wire      [3:0] src_pstrb,                                             // Write strobes
  output logic           src_pready,                                            // Ready
  output logic    [31:0] src_prdata,                                            // Read data
  // dst
  output logic     [9:0] dst_paddr,                                             // Address
  output logic           dst_psel,                                              // Select
  output logic           dst_penable,                                           // Enable
  output logic           dst_pwrite,                                            // Write not read
  output logic    [31:0] dst_pwdata,                                            // Write data
  output logic     [3:0] dst_pstrb,                                             // Write strobes
  input  wire            dst_pready,                                            // Ready
  input  wire     [31:0] dst_prdata                                             // Read data
);

logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (AXI4 subordinate)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Destination Port (AXI4 manager)
// ============================================
// Interface parameters
// APB Manager View
// APB Subordinate View
// APB Monitor View
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_apbtea5_epipe_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// Pipelining is disabled so feedthrough
assign dst_psel = src_psel;
assign dst_penable = src_penable;
assign dst_pwrite = src_pwrite;
assign dst_paddr = src_paddr;
assign dst_pwdata = src_pwdata;
assign dst_pstrb = src_pstrb;
assign src_pready = dst_pready;
assign src_prdata = dst_prdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_epipe_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea5_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea5_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea5_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_apbtea5_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_apbcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_wccg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_wdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_f1cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_rdcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_wdunpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wtr_req,
  output logic           wtr_rdy,
  input  wire      [2:0] wtr_size,                                              // Transfer size per data phase
  input  wire      [1:0] wtr_burst,                                             // Burst addressing mode
  input  wire     [11:0] wtr_addrlsb,                                           // 12 LSBs of address
  input  wire      [2:0] wtr_plen,                                              // Packet length in bytes
  output logic           w_valid,
  output logic    [31:0] w_data,
  output logic     [3:0] w_strb,
  output logic           w_last,
  input  wire            w_ready,
  input  wire            f_req,
  input  wire            f_eop,
  input  wire     [35:0] f_flitdata,
  output logic           f_ready,
  output logic    [11:0] wtr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [2:0] sizeCnvDiv;
logic     [4:0] firstCnt2Wrap;
logic     [7:0] wtr_mask;
logic     [7:0] wtr_mis;
logic    [10:0] firstXferCnt;
logic    [10:0] xferCnt;
logic    [10:0] xferCnt_nxt;
logic     [0:0] xferCnt_en;
logic    [10:0] useXferCnt;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic    [31:0] muxed_w_data;
logic     [3:0] muxed_w_strb;
logic           flitDone;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic     [0:0] haveFlit;
logic     [0:0] haveFlit_nxt;
logic     [0:0] haveFlit_en;
logic    [35:0] flitData;
logic    [35:0] flitData_nxt;
logic     [0:0] flitData_en;
logic           flitValid;
logic    [11:0] lower_baddr;
logic    [11:0] upper_baddr;
logic    [11:0] lower_addr;
logic    [11:0] upper_addr;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
logic    [11:0] saddr;
logic     [2:0] splen;
// Extracted from packet header
// APB W Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},wtr_plen} - 1'b1;                                    // We only care about 8 bits of address for our word indexing
assign wrapToAddr = wtr_addrlsb[7:0] & ~bamask;                                 // This is the address offset we wrap to
assign wrapIndex = wtr_addrlsb >> wtr_size;
assign sizeCnvDiv = wtr_plen >> wtr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign wtr_mask = (8'b1<<wtr_size) - 1'b1;
assign wtr_mis = wtr_addrlsb[7:0] & wtr_mask;
assign firstXferCnt = (wtr_burst!=2'd1) ? 11'(wtr_plen>>wtr_size) : 11'((16'(wtr_plen)+wtr_mask+wtr_mis)>>wtr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    xferCnt <= #1ps 11'd0;
  else if (xferCnt_en)
    xferCnt <= #1ps xferCnt_nxt;
end

assign useXferCnt = xferCnt;
always_comb
begin
  xferCnt_nxt = xferCnt;
  xferCnt_en  = 1'b0;
  if( newCmd )
    begin
      xferCnt_nxt = firstXferCnt;
      xferCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      xferCnt_nxt = useXferCnt - 1'd1;
      xferCnt_en  = 1'b1;
    end
end

assign wtr_rdy = ~trInPkt;
assign newCmd = wtr_req && wtr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = w_valid && w_ready;
assign f_ready = ~haveFlit || flitDone;
assign w_valid = flitValid;
assign w_last = w_valid && useXferCnt==11'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps wtr_burst;
end

assign use_tr_burst = held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps wtr_size;
end

assign use_tr_size = held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( busWriteValid && w_last )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> wtr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (wtr_addrlsb[7:0] & 8'd3) >> wtr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( w_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone;
assign muxed_w_data[7:0] = flitData[7:0];
assign muxed_w_strb[3:0] = flitData[35:32];
assign muxed_w_data[15:8] = flitData[15:8];
assign muxed_w_data[23:16] = flitData[23:16];
assign muxed_w_data[31:24] = flitData[31:24];
assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    haveFlit <= #1ps 1'd0;
  else if (haveFlit_en)
    haveFlit <= #1ps haveFlit_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitData <= #1ps {36{1'b0}};
  else if (flitData_en)
    flitData <= #1ps flitData_nxt;
end

assign flitValid = haveFlit;
always_comb
begin
  haveFlit_nxt   = haveFlit;
  haveFlit_en    = 1'b0;
  flitData_nxt   = flitData;
  flitData_en    = 1'b0;
  if( flitWriteValid )
    begin
      haveFlit_nxt   = 1'b1;
      haveFlit_en    = 1'b1;
      flitData_en    = 1'b1;
      flitData_nxt   = f_flitdata;
    end
  else if( flitDone )
    begin
      haveFlit_nxt   = 1'b0;
      haveFlit_en    = 1'b1;
    end
end

assign w_data[7:0] = (w_valid && wrMask[0]) ? muxed_w_data[7:0] : 8'd0;
assign w_data[15:8] = (w_valid && wrMask[1]) ? muxed_w_data[15:8] : 8'd0;
assign w_data[23:16] = (w_valid && wrMask[2]) ? muxed_w_data[23:16] : 8'd0;
assign w_data[31:24] = (w_valid && wrMask[3]) ? muxed_w_data[31:24] : 8'd0;
assign w_strb = w_valid ? muxed_w_strb & wrMask : 4'd0;
assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  addrlsb_nxt   = addrlsb;
  // Write enables
  addrlsb_en    = 1'b0;
  if (newCmd)
    begin
      addrlsb_nxt = wtr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred from packing FIFO
  else if (busWriteValid)
    begin
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps wtr_addrlsb;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps wtr_plen;
end

assign wtr_addrlsb_out = !(newCmd) ? addrlsb : wtr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_apbtea5_rdpack (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            tr_req,
  output logic           tr_rdy,
  input  wire      [2:0] tr_size,
  input  wire      [1:0] tr_burst,
  input  wire     [11:0] tr_addrlsb,
  input  wire      [2:0] tr_plen,
  output logic           r_req,
  output logic           r_last,
  input  wire     [31:0] r_data,
  input  wire            r_slverr,
  input  wire            r_ready,
  output logic           f_req,
  output logic           f_eop,
  output logic    [33:0] f_flitdata,
  input  wire            f_ready,
  output logic    [11:0] tr_addrlsb_out
);

logic     [7:0] bamask;                                                         // We only care about 8 bits of address for our word indexing
logic     [7:0] wrapToAddr;                                                     // This is the address offset we wrap to
logic    [11:0] wrapIndex;
logic     [4:0] firstCnt2Wrap;
logic     [2:0] sizeCnvDiv;
logic           newCmd;
logic           flitWriteValid;
logic           busWriteValid;
logic     [0:0] heldFlitDone;
logic     [0:0] heldEop;
logic     [1:0] held_tr_burst;
logic     [1:0] use_tr_burst;
logic     [2:0] held_tr_size;
logic     [2:0] use_tr_size;
logic           isFixed;
logic           isNarrow;
logic           isWrap;
logic     [0:0] trInPkt;
logic     [0:0] trInPkt_nxt;
logic     [0:0] trInPkt_en;
logic     [7:0] subBusWdCntWrap_tmp;
logic     [1:0] subBusWdCntWrap;
logic     [1:0] subBusWdCntWrap_nxt;
logic     [1:0] useSubBusWdCntWrap;
logic     [4:0] cnt2Wrap;
logic     [4:0] cnt2Wrap_nxt;
logic     [0:0] cnt2Wrap_en;
logic     [4:0] useCnt2Wrap;
logic           busWdWrap;
logic     [7:0] firstSubBusWdCnt;
logic     [7:0] subBusWdMax;
logic     [1:0] subBusWdCnt;
logic     [1:0] subBusWdCnt_nxt;
logic     [0:0] subBusWdCnt_en;
logic     [1:0] useSubBusWdCnt;
logic           busWdDone;
logic           flitDone;
logic           useBusWdCnt;
logic    [33:0] flitWd;
logic    [33:0] flitWd_nxt;
logic     [0:0] flitWd_en;
logic     [7:0] size;
logic     [7:0] unused;
logic     [3:0] preMask;
logic     [3:0] wrMask;
logic    [11:0] esize;
logic    [11:0] amask;
logic    [11:0] bamask12;                                                       // Burst address mask is transfer length minus 1 // 
logic    [11:0] lower_baddr;                                                    // Lower burst address
logic    [11:0] upper_baddr;                                                    // Upper burst address
logic    [11:0] lower_addr;                                                     // Lower element address
logic    [11:0] upper_addr;                                                     // Upper element address
logic    [11:0] esize_minus_first_offset;
logic    [11:0] first_offset;
logic     [2:0] raw_wcnt;
logic     [2:0] wcnt;
logic    [11:0] saddr;
logic     [2:0] wplen;
logic     [2:0] wplen_nxt;
logic     [0:0] wplen_en;
logic     [2:0] splen;
logic    [11:0] addrlsb;
logic    [11:0] addrlsb_nxt;
logic     [0:0] addrlsb_en;
// Extracted from AXI AW Channel
// APB R Channel
// Flit Bus
// Incrementing address
assign bamask = {{5{1'b0}},tr_plen} - 1'b1;                                     // We only care about 8 bits of address for our word indexing
assign wrapToAddr = tr_addrlsb[7:0] & ~bamask;                                  // This is the address offset we wrap to
assign wrapIndex = tr_addrlsb >> tr_size;
assign firstCnt2Wrap = {{2{1'b0}},sizeCnvDiv} - (wrapIndex[4:0] & ({{2{1'b0}},sizeCnvDiv}-5'b1));
assign sizeCnvDiv = tr_plen >> tr_size;
assign tr_rdy = ~trInPkt;
assign f_flitdata = flitWd;
assign f_req = heldFlitDone;
assign f_eop = heldEop;
assign r_req = trInPkt_nxt && (!heldFlitDone || flitWriteValid);
assign newCmd = tr_req && tr_rdy;
assign flitWriteValid = f_req && f_ready;
assign busWriteValid = r_ready && r_req;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldFlitDone <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldFlitDone <= #1ps flitDone;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    heldEop <= #1ps 1'd0;
  else if (flitDone || flitWriteValid)
    heldEop <= #1ps flitDone && r_last;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_burst <= #1ps 2'd0;
  else if (newCmd)
    held_tr_burst <= #1ps tr_burst;
end

assign use_tr_burst = (newCmd) ? tr_burst : held_tr_burst;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    held_tr_size <= #1ps 3'd0;
  else if (newCmd)
    held_tr_size <= #1ps tr_size;
end

assign use_tr_size = (newCmd) ? tr_size : held_tr_size;
assign isFixed = (use_tr_burst==2'd0);
assign isNarrow = use_tr_size<3'd2;
assign isWrap = (use_tr_burst==2'd2);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    trInPkt <= #1ps 1'd0;
  else if (trInPkt_en)
    trInPkt <= #1ps trInPkt_nxt;
end

always_comb
begin
  trInPkt_nxt = trInPkt;
  trInPkt_en  = 1'b0;
  if( newCmd )
    begin
      trInPkt_nxt = 1'b1;
      trInPkt_en  = 1'b1;
    end
  if( flitWriteValid && f_eop )
    begin
      trInPkt_nxt = 1'b0;
      trInPkt_en  = 1'b1;
    end
end

assign subBusWdCntWrap_tmp = (wrapToAddr & 8'd3) >> tr_size;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCntWrap <= #1ps 2'd0;
  else if (newCmd)
    subBusWdCntWrap <= #1ps subBusWdCntWrap_nxt;
end

assign subBusWdCntWrap_nxt = subBusWdCntWrap_tmp[1:0];
assign useSubBusWdCntWrap = (newCmd) ? subBusWdCntWrap_nxt : subBusWdCntWrap;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    cnt2Wrap <= #1ps 5'd0;
  else if (cnt2Wrap_en)
    cnt2Wrap <= #1ps cnt2Wrap_nxt;
end

assign useCnt2Wrap = newCmd ? firstCnt2Wrap : cnt2Wrap;
always_comb
begin
  cnt2Wrap_nxt = cnt2Wrap;
  cnt2Wrap_en  = 1'b0;
  busWdWrap    = 1'b0;
  if(newCmd)
    begin
      cnt2Wrap_nxt = firstCnt2Wrap;
      cnt2Wrap_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      cnt2Wrap_nxt = useCnt2Wrap - 5'd1;
      cnt2Wrap_en  = 1'b1;
      if( useCnt2Wrap==5'd1 )
        begin
          busWdWrap = isWrap;
        end
    end
end

assign firstSubBusWdCnt = (tr_addrlsb[7:0] & 8'd3) >> tr_size;
assign subBusWdMax = (8'd4 >> use_tr_size) - 8'd1;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    subBusWdCnt <= #1ps 2'd0;
  else if (subBusWdCnt_en)
    subBusWdCnt <= #1ps subBusWdCnt_nxt;
end

assign useSubBusWdCnt = (newCmd) ? firstSubBusWdCnt[1:0] : subBusWdCnt;
always_comb
begin
  subBusWdCnt_nxt = subBusWdCnt;
  subBusWdCnt_en  = 1'b0;
  busWdDone       = 1'b0;
  if( newCmd )
    begin
      subBusWdCnt_nxt = firstSubBusWdCnt[1:0];
      subBusWdCnt_en  = 1'b1;
    end
  if( busWriteValid )
    begin
      if( r_last || isFixed )
          busWdDone = 1'b1;
      else if( busWdWrap )
        begin
          subBusWdCnt_nxt = useSubBusWdCntWrap;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else if( useSubBusWdCnt == subBusWdMax[1:0] )
        begin
          subBusWdCnt_nxt = 2'd0;
          subBusWdCnt_en  = 1'b1;
          busWdDone = 1'b1;
        end
      else
        begin
          subBusWdCnt_nxt = useSubBusWdCnt + 2'd1;
          subBusWdCnt_en  = 1'b1;
        end
    end
end

assign flitDone = busWdDone || (isNarrow && busWriteValid);
assign useBusWdCnt = 1'b0;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    flitWd <= #1ps {34{1'b0}};
  else if (flitWd_en)
    flitWd <= #1ps flitWd_nxt;
end

assign size = (8'd1<<use_tr_size);
assign unused = 8'd4 - size;
assign preMask = {4{1'b1}} >> unused;
assign wrMask = preMask << ({{5{1'b0}},useSubBusWdCnt}<<use_tr_size);
always_comb
begin
  // First, assign the bus word to every possible flit word slot
  flitWd_nxt = flitWriteValid ? {34{1'b0}} : flitWd;
  // Start out with nothing enabled
  flitWd_en = flitWriteValid ? 1'b1 : 1'b0;
  // Now enable any bytes that are being written this cycle
  if( busWriteValid )
    begin
      if( useBusWdCnt == 1'd0 )
        begin
          if( wrMask[0] )
            begin
              flitWd_nxt[7:0] = r_data[7:0];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[1] )
            begin
              flitWd_nxt[15:8] = r_data[15:8];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[2] )
            begin
              flitWd_nxt[23:16] = r_data[23:16];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
          if( wrMask[3] )
            begin
              flitWd_nxt[31:24] = r_data[31:24];
              flitWd_nxt[33:32] = {r_slverr, 1'b0};
              flitWd_en         = 1'b1;
            end
        end
    end
end

assign esize = 12'd1 << use_tr_size;
assign amask = esize - 12'd1;
assign bamask12 = {{9{1'b0}},splen} - 1'b1;                                     // Burst address mask is transfer length minus 1 // 
assign lower_baddr = saddr & ~bamask12;                                         // Lower burst address
assign upper_baddr = lower_baddr + {{9{1'b0}},splen};                           // Upper burst address
assign lower_addr = addrlsb & ~amask;                                           // Lower element address
assign upper_addr = lower_addr + esize;                                         // Upper element address
assign esize_minus_first_offset = esize - first_offset;
assign first_offset = addrlsb & amask;
assign raw_wcnt = (held_tr_burst == 2'd1) ? esize_minus_first_offset[2:0] : esize[2:0];
assign wcnt = (raw_wcnt > wplen) ? wplen : raw_wcnt;
assign r_last = (wcnt >= wplen);
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    saddr <= #1ps 12'd0;
  else if (newCmd)
    saddr <= #1ps tr_addrlsb;
end

// Write remaining packet length and address LSB tracking flops
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    wplen <= #1ps 3'd0;
  else if (wplen_en)
    wplen <= #1ps wplen_nxt;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    splen <= #1ps 3'd0;
  else if (newCmd)
    splen <= #1ps tr_plen;
end

always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    addrlsb <= #1ps 12'd0;
  else if (addrlsb_en)
    addrlsb <= #1ps addrlsb_nxt;
end

// Write Address and count tracking
always_comb
begin
  // Defaults
  wplen_nxt   = wplen;
  addrlsb_nxt = addrlsb;
  wplen_en    = 1'b0;
  addrlsb_en  = 1'b0;
  if (tr_req && tr_rdy)
    begin
      wplen_nxt   = tr_plen;
      wplen_en    = 1'b1;
      addrlsb_nxt = tr_addrlsb;
      addrlsb_en  = 1'b1;
    end
  // Data was transferred to packing FIFO
  else if (busWriteValid)
    begin
      wplen_en    = 1'b1;
      addrlsb_en  = 1'b1;
      // Generate next address LSBs (and input byte positions)
      case (held_tr_burst)
        // Fixed Burst
        2'd0:
          begin
            wplen_nxt   = wplen - wcnt;
            addrlsb_nxt = addrlsb;
          end
        // Linear Incrementing
        2'd1:
          begin
            wplen_nxt   = wplen   - wcnt;
            addrlsb_nxt = upper_addr;
          end
        // Wrap
        2'd2:
          begin
            wplen_nxt   = wplen      - wcnt;
            if (upper_addr == upper_baddr)
              addrlsb_nxt = lower_baddr;
            else
              addrlsb_nxt = upper_addr;
          end
        default:
          begin
            wplen_nxt   = wplen;
            addrlsb_nxt = upper_addr;
          end
      endcase
    end
end

assign tr_addrlsb_out = !(newCmd) ? addrlsb : tr_addrlsb;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0 (
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  // slf0
  input  wire            slf0_activity,                                         // Upcoming activity indicator
  input  wire            slf0_req,                                              // Flit transfer request
  input  wire            slf0_sop,                                              // Start of packet indicator
  input  wire            slf0_eop,                                              // End of packet indicator
  input  wire     [35:0] slf0_flitdata,                                         // Flit data
  output logic           slf0_ready,                                            // Flit transfer ready
  // slf1
  input  wire            slf1_activity,                                         // Upcoming activity indicator
  input  wire            slf1_req,                                              // Flit transfer request
  input  wire            slf1_sop,                                              // Start of packet indicator
  input  wire            slf1_eop,                                              // End of packet indicator
  input  wire     [59:0] slf1_flitdata,                                         // Flit data
  output logic           slf1_ready,                                            // Flit transfer ready
  // slr0
  output logic           slr0_activity,                                         // Upcoming activity indicator
  output logic           slr0_req,                                              // Flit transfer request
  output logic           slr0_sop,                                              // Start of packet indicator
  output logic           slr0_eop,                                              // End of packet indicator
  output logic    [33:0] slr0_flitdata,                                         // Flit data
  input  wire            slr0_ready,                                            // Flit transfer ready
  // slr1
  output logic           slr1_activity,                                         // Upcoming activity indicator
  output logic           slr1_req,                                              // Flit transfer request
  output logic           slr1_sop,                                              // Start of packet indicator
  output logic           slr1_eop,                                              // End of packet indicator
  output logic    [23:0] slr1_flitdata,                                         // Flit data
  input  wire            slr1_ready,                                            // Flit transfer ready
  // dlf0
  output logic           dlf0_activity,                                         // Upcoming activity indicator
  output logic           dlf0_req,                                              // Flit transfer request
  output logic           dlf0_sop,                                              // Start of packet indicator
  output logic           dlf0_eop,                                              // End of packet indicator
  output logic    [35:0] dlf0_flitdata,                                         // Flit data
  input  wire            dlf0_ready,                                            // Flit transfer ready
  // dlf1
  output logic           dlf1_activity,                                         // Upcoming activity indicator
  output logic           dlf1_req,                                              // Flit transfer request
  output logic           dlf1_sop,                                              // Start of packet indicator
  output logic           dlf1_eop,                                              // End of packet indicator
  output logic    [59:0] dlf1_flitdata,                                         // Flit data
  input  wire            dlf1_ready,                                            // Flit transfer ready
  // dlr0
  input  wire            dlr0_activity,                                         // Upcoming activity indicator
  input  wire            dlr0_req,                                              // Flit transfer request
  input  wire            dlr0_sop,                                              // Start of packet indicator
  input  wire            dlr0_eop,                                              // End of packet indicator
  input  wire     [33:0] dlr0_flitdata,                                         // Flit data
  output logic           dlr0_ready,                                            // Flit transfer ready
  // dlr1
  input  wire            dlr1_activity,                                         // Upcoming activity indicator
  input  wire            dlr1_req,                                              // Flit transfer request
  input  wire            dlr1_sop,                                              // Start of packet indicator
  input  wire            dlr1_eop,                                              // End of packet indicator
  input  wire     [23:0] dlr1_flitdata,                                         // Flit data
  output logic           dlr1_ready                                             // Flit transfer ready
);

logic           glk_f0_0_activity;                                              // Upcoming activity indicator
logic           glk_f0_0_strb;                                                  // Flit transfer strobe
logic           glk_f0_0_sop;                                                   // Start of Packet Flit Indicator
logic           glk_f0_0_eop;                                                   // End of Packet Flit Indicator
logic    [35:0] glk_f0_0_flitdata;                                              // Flit data
logic           glk_f0_0_ret_activity;                                          // Upcoming credit return activity indicator
logic           glk_f0_0_ret_strb;                                              // Credit return strobe
logic     [0:0] glk_f0_0_ret_cnt;                                               // Credit return credit count
logic           glk_f1_0_activity;                                              // Upcoming activity indicator
logic           glk_f1_0_strb;                                                  // Flit transfer strobe
logic           glk_f1_0_sop;                                                   // Start of Packet Flit Indicator
logic           glk_f1_0_eop;                                                   // End of Packet Flit Indicator
logic    [59:0] glk_f1_0_flitdata;                                              // Flit data
logic           glk_f1_0_ret_activity;                                          // Upcoming credit return activity indicator
logic           glk_f1_0_ret_strb;                                              // Credit return strobe
logic     [0:0] glk_f1_0_ret_cnt;                                               // Credit return credit count
logic           glk_r0_0_activity;                                              // Upcoming activity indicator
logic           glk_r0_0_strb;                                                  // Flit transfer strobe
logic           glk_r0_0_sop;                                                   // Start of Packet Flit Indicator
logic           glk_r0_0_eop;                                                   // End of Packet Flit Indicator
logic    [33:0] glk_r0_0_flitdata;                                              // Flit data
logic           glk_r0_0_ret_activity;                                          // Upcoming credit return activity indicator
logic           glk_r0_0_ret_strb;                                              // Credit return strobe
logic     [0:0] glk_r0_0_ret_cnt;                                               // Credit return credit count
logic           glk_r1_0_activity;                                              // Upcoming activity indicator
logic           glk_r1_0_strb;                                                  // Flit transfer strobe
logic           glk_r1_0_sop;                                                   // Start of Packet Flit Indicator
logic           glk_r1_0_eop;                                                   // End of Packet Flit Indicator
logic    [23:0] glk_r1_0_flitdata;                                              // Flit data
logic           glk_r1_0_ret_activity;                                          // Upcoming credit return activity indicator
logic           glk_r1_0_ret_strb;                                              // Credit return strobe
logic     [0:0] glk_r1_0_ret_cnt;                                               // Credit return credit count
// Source clock / reset (may be only)
// Destination clock / reset (may be only)
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Side LLK Forward Channels (LLK manager)
// ============================================
// ============================================
// Source Side LLK Reverse Channels (LLK subordinate)
// ============================================
// ============================================
// Dest Side LLK Forward Channels (LLK manager)
// ============================================
// ============================================
// Dest Side LLK Reverse Channels (LLK subordinate)
// ============================================
// ===========================================
// NoC Link Source Instance
// ===========================================
usb4_tc_noc_link0_ls ls (
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .llk_f0_activity(slf0_activity),                                              // i:1
  .llk_f0_req(slf0_req),                                                        // i:1
  .llk_f0_sop(slf0_sop),                                                        // i:1
  .llk_f0_eop(slf0_eop),                                                        // i:1
  .llk_f0_flitdata(slf0_flitdata),                                              // i:36
  .llk_f0_ready(slf0_ready),                                                    // o:1
  .llk_f1_activity(slf1_activity),                                              // i:1
  .llk_f1_req(slf1_req),                                                        // i:1
  .llk_f1_sop(slf1_sop),                                                        // i:1
  .llk_f1_eop(slf1_eop),                                                        // i:1
  .llk_f1_flitdata(slf1_flitdata),                                              // i:60
  .llk_f1_ready(slf1_ready),                                                    // o:1
  .llk_r0_activity(slr0_activity),                                              // o:1
  .llk_r0_req(slr0_req),                                                        // o:1
  .llk_r0_sop(slr0_sop),                                                        // o:1
  .llk_r0_eop(slr0_eop),                                                        // o:1
  .llk_r0_flitdata(slr0_flitdata),                                              // o:34
  .llk_r0_ready(slr0_ready),                                                    // i:1
  .llk_r1_activity(slr1_activity),                                              // o:1
  .llk_r1_req(slr1_req),                                                        // o:1
  .llk_r1_sop(slr1_sop),                                                        // o:1
  .llk_r1_eop(slr1_eop),                                                        // o:1
  .llk_r1_flitdata(slr1_flitdata),                                              // o:24
  .llk_r1_ready(slr1_ready),                                                    // i:1
  .glk_f0_activity(glk_f0_0_activity),                                          // o:1
  .glk_f0_strb(glk_f0_0_strb),                                                  // o:1
  .glk_f0_sop(glk_f0_0_sop),                                                    // o:1
  .glk_f0_eop(glk_f0_0_eop),                                                    // o:1
  .glk_f0_flitdata(glk_f0_0_flitdata),                                          // o:36
  .glk_f0_ret_activity(glk_f0_0_ret_activity),                                  // i:1
  .glk_f0_ret_strb(glk_f0_0_ret_strb),                                          // i:1
  .glk_f0_ret_cnt(glk_f0_0_ret_cnt),                                            // i:1
  .glk_f1_activity(glk_f1_0_activity),                                          // o:1
  .glk_f1_strb(glk_f1_0_strb),                                                  // o:1
  .glk_f1_sop(glk_f1_0_sop),                                                    // o:1
  .glk_f1_eop(glk_f1_0_eop),                                                    // o:1
  .glk_f1_flitdata(glk_f1_0_flitdata),                                          // o:60
  .glk_f1_ret_activity(glk_f1_0_ret_activity),                                  // i:1
  .glk_f1_ret_strb(glk_f1_0_ret_strb),                                          // i:1
  .glk_f1_ret_cnt(glk_f1_0_ret_cnt),                                            // i:1
  .glk_r0_activity(glk_r0_0_activity),                                          // i:1
  .glk_r0_strb(glk_r0_0_strb),                                                  // i:1
  .glk_r0_sop(glk_r0_0_sop),                                                    // i:1
  .glk_r0_eop(glk_r0_0_eop),                                                    // i:1
  .glk_r0_flitdata(glk_r0_0_flitdata),                                          // i:34
  .glk_r0_ret_activity(glk_r0_0_ret_activity),                                  // o:1
  .glk_r0_ret_strb(glk_r0_0_ret_strb),                                          // o:1
  .glk_r0_ret_cnt(glk_r0_0_ret_cnt),                                            // o:1
  .glk_r1_activity(glk_r1_0_activity),                                          // i:1
  .glk_r1_strb(glk_r1_0_strb),                                                  // i:1
  .glk_r1_sop(glk_r1_0_sop),                                                    // i:1
  .glk_r1_eop(glk_r1_0_eop),                                                    // i:1
  .glk_r1_flitdata(glk_r1_0_flitdata),                                          // i:24
  .glk_r1_ret_activity(glk_r1_0_ret_activity),                                  // o:1
  .glk_r1_ret_strb(glk_r1_0_ret_strb),                                          // o:1
  .glk_r1_ret_cnt(glk_r1_0_ret_cnt)                                             // o:1
);
// ===========================================
// NoC Link Target Instance
// ===========================================
usb4_tc_noc_link0_lt lt (
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .glk_f0_activity(glk_f0_0_activity),                                          // i:1
  .glk_f0_strb(glk_f0_0_strb),                                                  // i:1
  .glk_f0_sop(glk_f0_0_sop),                                                    // i:1
  .glk_f0_eop(glk_f0_0_eop),                                                    // i:1
  .glk_f0_flitdata(glk_f0_0_flitdata),                                          // i:36
  .glk_f0_ret_activity(glk_f0_0_ret_activity),                                  // o:1
  .glk_f0_ret_strb(glk_f0_0_ret_strb),                                          // o:1
  .glk_f0_ret_cnt(glk_f0_0_ret_cnt),                                            // o:1
  .glk_f1_activity(glk_f1_0_activity),                                          // i:1
  .glk_f1_strb(glk_f1_0_strb),                                                  // i:1
  .glk_f1_sop(glk_f1_0_sop),                                                    // i:1
  .glk_f1_eop(glk_f1_0_eop),                                                    // i:1
  .glk_f1_flitdata(glk_f1_0_flitdata),                                          // i:60
  .glk_f1_ret_activity(glk_f1_0_ret_activity),                                  // o:1
  .glk_f1_ret_strb(glk_f1_0_ret_strb),                                          // o:1
  .glk_f1_ret_cnt(glk_f1_0_ret_cnt),                                            // o:1
  .glk_r0_activity(glk_r0_0_activity),                                          // o:1
  .glk_r0_strb(glk_r0_0_strb),                                                  // o:1
  .glk_r0_sop(glk_r0_0_sop),                                                    // o:1
  .glk_r0_eop(glk_r0_0_eop),                                                    // o:1
  .glk_r0_flitdata(glk_r0_0_flitdata),                                          // o:34
  .glk_r0_ret_activity(glk_r0_0_ret_activity),                                  // i:1
  .glk_r0_ret_strb(glk_r0_0_ret_strb),                                          // i:1
  .glk_r0_ret_cnt(glk_r0_0_ret_cnt),                                            // i:1
  .glk_r1_activity(glk_r1_0_activity),                                          // o:1
  .glk_r1_strb(glk_r1_0_strb),                                                  // o:1
  .glk_r1_sop(glk_r1_0_sop),                                                    // o:1
  .glk_r1_eop(glk_r1_0_eop),                                                    // o:1
  .glk_r1_flitdata(glk_r1_0_flitdata),                                          // o:24
  .glk_r1_ret_activity(glk_r1_0_ret_activity),                                  // i:1
  .glk_r1_ret_strb(glk_r1_0_ret_strb),                                          // i:1
  .glk_r1_ret_cnt(glk_r1_0_ret_cnt),                                            // i:1
  .llk_f0_activity(dlf0_activity),                                              // o:1
  .llk_f0_req(dlf0_req),                                                        // o:1
  .llk_f0_sop(dlf0_sop),                                                        // o:1
  .llk_f0_eop(dlf0_eop),                                                        // o:1
  .llk_f0_flitdata(dlf0_flitdata),                                              // o:36
  .llk_f0_ready(dlf0_ready),                                                    // i:1
  .llk_f1_activity(dlf1_activity),                                              // o:1
  .llk_f1_req(dlf1_req),                                                        // o:1
  .llk_f1_sop(dlf1_sop),                                                        // o:1
  .llk_f1_eop(dlf1_eop),                                                        // o:1
  .llk_f1_flitdata(dlf1_flitdata),                                              // o:60
  .llk_f1_ready(dlf1_ready),                                                    // i:1
  .llk_r0_activity(dlr0_activity),                                              // i:1
  .llk_r0_req(dlr0_req),                                                        // i:1
  .llk_r0_sop(dlr0_sop),                                                        // i:1
  .llk_r0_eop(dlr0_eop),                                                        // i:1
  .llk_r0_flitdata(dlr0_flitdata),                                              // i:34
  .llk_r0_ready(dlr0_ready),                                                    // o:1
  .llk_r1_activity(dlr1_activity),                                              // i:1
  .llk_r1_req(dlr1_req),                                                        // i:1
  .llk_r1_sop(dlr1_sop),                                                        // i:1
  .llk_r1_eop(dlr1_eop),                                                        // i:1
  .llk_r1_flitdata(dlr1_flitdata),                                              // i:24
  .llk_r1_ready(dlr1_ready)                                                     // o:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls (
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  // llk_f0
  input  wire            llk_f0_activity,                                       // Upcoming activity indicator
  input  wire            llk_f0_req,                                            // Flit transfer request
  input  wire            llk_f0_sop,                                            // Start of packet indicator
  input  wire            llk_f0_eop,                                            // End of packet indicator
  input  wire     [35:0] llk_f0_flitdata,                                       // Flit data
  output logic           llk_f0_ready,                                          // Flit transfer ready
  // llk_f1
  input  wire            llk_f1_activity,                                       // Upcoming activity indicator
  input  wire            llk_f1_req,                                            // Flit transfer request
  input  wire            llk_f1_sop,                                            // Start of packet indicator
  input  wire            llk_f1_eop,                                            // End of packet indicator
  input  wire     [59:0] llk_f1_flitdata,                                       // Flit data
  output logic           llk_f1_ready,                                          // Flit transfer ready
  // llk_r0
  output logic           llk_r0_activity,                                       // Upcoming activity indicator
  output logic           llk_r0_req,                                            // Flit transfer request
  output logic           llk_r0_sop,                                            // Start of packet indicator
  output logic           llk_r0_eop,                                            // End of packet indicator
  output logic    [33:0] llk_r0_flitdata,                                       // Flit data
  input  wire            llk_r0_ready,                                          // Flit transfer ready
  // llk_r1
  output logic           llk_r1_activity,                                       // Upcoming activity indicator
  output logic           llk_r1_req,                                            // Flit transfer request
  output logic           llk_r1_sop,                                            // Start of packet indicator
  output logic           llk_r1_eop,                                            // End of packet indicator
  output logic    [23:0] llk_r1_flitdata,                                       // Flit data
  input  wire            llk_r1_ready,                                          // Flit transfer ready
  // glk_f0
  output logic           glk_f0_activity,                                       // Upcoming activity indicator
  output logic           glk_f0_strb,                                           // Flit transfer strobe
  output logic           glk_f0_sop,                                            // Start of Packet Flit Indicator
  output logic           glk_f0_eop,                                            // End of Packet Flit Indicator
  output logic    [35:0] glk_f0_flitdata,                                       // Flit data
  input  wire            glk_f0_ret_activity,                                   // Upcoming credit return activity indicator
  input  wire            glk_f0_ret_strb,                                       // Credit return strobe
  input  wire      [0:0] glk_f0_ret_cnt,                                        // Credit return credit count
  // glk_f1
  output logic           glk_f1_activity,                                       // Upcoming activity indicator
  output logic           glk_f1_strb,                                           // Flit transfer strobe
  output logic           glk_f1_sop,                                            // Start of Packet Flit Indicator
  output logic           glk_f1_eop,                                            // End of Packet Flit Indicator
  output logic    [59:0] glk_f1_flitdata,                                       // Flit data
  input  wire            glk_f1_ret_activity,                                   // Upcoming credit return activity indicator
  input  wire            glk_f1_ret_strb,                                       // Credit return strobe
  input  wire      [0:0] glk_f1_ret_cnt,                                        // Credit return credit count
  // glk_r0
  input  wire            glk_r0_activity,                                       // Upcomong activity indicator
  input  wire            glk_r0_strb,                                           // Request
  input  wire            glk_r0_sop,                                            // Start of Packet Flit Indicator
  input  wire            glk_r0_eop,                                            // End of Packet Flit Indicator
  input  wire     [33:0] glk_r0_flitdata,                                       // Flit data
  output logic           glk_r0_ret_activity,                                   // Upcoming credit return activity indicator
  output logic           glk_r0_ret_strb,                                       // Credit return strobe
  output logic     [0:0] glk_r0_ret_cnt,                                        // Credit return credit count
  // glk_r1
  input  wire            glk_r1_activity,                                       // Upcomong activity indicator
  input  wire            glk_r1_strb,                                           // Request
  input  wire            glk_r1_sop,                                            // Start of Packet Flit Indicator
  input  wire            glk_r1_eop,                                            // End of Packet Flit Indicator
  input  wire     [23:0] glk_r1_flitdata,                                       // Flit data
  output logic           glk_r1_ret_activity,                                   // Upcoming credit return activity indicator
  output logic           glk_r1_ret_strb,                                       // Credit return strobe
  output logic     [0:0] glk_r1_ret_cnt                                         // Credit return credit count
);

// =========================================================
// Clocks / Resets
// =========================================================
// Local clock / reset (may be only clock / reset)
// Global clock / reset
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// =========================================================
// Source Side LLK Forward Channel Interfces (LLK manager)
// =========================================================
// =========================================================
// LLK Reverse Channel Interfaces (LLK subordinate)
// =========================================================
// =========================================================
// LK Forward Channel Interfaces (LK manager)
// =========================================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// =========================================================
// LK Reverse Channel Interfaces (LK subordinate)
// =========================================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// NoC L2G Bridge Instances
// ===========================================
usb4_tc_noc_link0_ls_l2g_f0 l2g_f0 (
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .llk_activity(llk_f0_activity),                                               // i:1
  .llk_req(llk_f0_req),                                                         // i:1
  .llk_sop(llk_f0_sop),                                                         // i:1
  .llk_eop(llk_f0_eop),                                                         // i:1
  .llk_flitdata(llk_f0_flitdata),                                               // i:36
  .llk_ready(llk_f0_ready),                                                     // o:1
  .glk_activity(glk_f0_activity),                                               // o:1
  .glk_strb(glk_f0_strb),                                                       // o:1
  .glk_sop(glk_f0_sop),                                                         // o:1
  .glk_eop(glk_f0_eop),                                                         // o:1
  .glk_flitdata(glk_f0_flitdata),                                               // o:36
  .glk_ret_activity(glk_f0_ret_activity),                                       // i:1
  .glk_ret_strb(glk_f0_ret_strb),                                               // i:1
  .glk_ret_cnt(glk_f0_ret_cnt)                                                  // i:1
);
usb4_tc_noc_link0_ls_l2g_f1 l2g_f1 (
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .llk_activity(llk_f1_activity),                                               // i:1
  .llk_req(llk_f1_req),                                                         // i:1
  .llk_sop(llk_f1_sop),                                                         // i:1
  .llk_eop(llk_f1_eop),                                                         // i:1
  .llk_flitdata(llk_f1_flitdata),                                               // i:60
  .llk_ready(llk_f1_ready),                                                     // o:1
  .glk_activity(glk_f1_activity),                                               // o:1
  .glk_strb(glk_f1_strb),                                                       // o:1
  .glk_sop(glk_f1_sop),                                                         // o:1
  .glk_eop(glk_f1_eop),                                                         // o:1
  .glk_flitdata(glk_f1_flitdata),                                               // o:60
  .glk_ret_activity(glk_f1_ret_activity),                                       // i:1
  .glk_ret_strb(glk_f1_ret_strb),                                               // i:1
  .glk_ret_cnt(glk_f1_ret_cnt)                                                  // i:1
);
// ===========================================
// NoC G2L Bridge Instances
// ===========================================
usb4_tc_noc_link0_ls_g2l_r0 g2l_r0 (
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .glk_activity(glk_r0_activity),                                               // i:1
  .glk_strb(glk_r0_strb),                                                       // i:1
  .glk_sop(glk_r0_sop),                                                         // i:1
  .glk_eop(glk_r0_eop),                                                         // i:1
  .glk_flitdata(glk_r0_flitdata),                                               // i:34
  .glk_ret_activity(glk_r0_ret_activity),                                       // o:1
  .glk_ret_strb(glk_r0_ret_strb),                                               // o:1
  .glk_ret_cnt(glk_r0_ret_cnt),                                                 // o:1
  .llk_activity(llk_r0_activity),                                               // o:1
  .llk_req(llk_r0_req),                                                         // o:1
  .llk_sop(llk_r0_sop),                                                         // o:1
  .llk_eop(llk_r0_eop),                                                         // o:1
  .llk_flitdata(llk_r0_flitdata),                                               // o:34
  .llk_ready(llk_r0_ready)                                                      // i:1
);
usb4_tc_noc_link0_ls_g2l_r1 g2l_r1 (
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .glk_activity(glk_r1_activity),                                               // i:1
  .glk_strb(glk_r1_strb),                                                       // i:1
  .glk_sop(glk_r1_sop),                                                         // i:1
  .glk_eop(glk_r1_eop),                                                         // i:1
  .glk_flitdata(glk_r1_flitdata),                                               // i:24
  .glk_ret_activity(glk_r1_ret_activity),                                       // o:1
  .glk_ret_strb(glk_r1_ret_strb),                                               // o:1
  .glk_ret_cnt(glk_r1_ret_cnt),                                                 // o:1
  .llk_activity(llk_r1_activity),                                               // o:1
  .llk_req(llk_r1_req),                                                         // o:1
  .llk_sop(llk_r1_sop),                                                         // o:1
  .llk_eop(llk_r1_eop),                                                         // o:1
  .llk_flitdata(llk_r1_flitdata),                                               // o:24
  .llk_ready(llk_r1_ready)                                                      // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f0 (
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  // llk
  input  wire            llk_activity,                                          // Upcoming activity indicator
  input  wire            llk_req,                                               // Flit transfer request
  input  wire            llk_sop,                                               // Start of packet indicator
  input  wire            llk_eop,                                               // End of packet indicator
  input  wire     [35:0] llk_flitdata,                                          // Flit data
  output logic           llk_ready,                                             // Flit transfer ready
  // glk
  output logic           glk_activity,                                          // Upcoming activity indicator
  output logic           glk_strb,                                              // Flit transfer strobe
  output logic           glk_sop,                                               // Start of Packet Flit Indicator
  output logic           glk_eop,                                               // End of Packet Flit Indicator
  output logic    [35:0] glk_flitdata,                                          // Flit data
  input  wire            glk_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            glk_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] glk_ret_cnt                                            // Credit return credit count
);

logic           glkp_activity;                                                  // Upcomong activity indicator
logic           glkp_strb;                                                      // Request
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [35:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [35:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           credclk;
logic           credclkAct;
wire            credclkEn;
logic    [11:0] ccnt;
logic    [11:0] ccnt_nxt;
logic     [0:0] ccnt_en;
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// LLK Interface
// ============================================
// ============================================
// LK Interface
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_l2g_f0_gpipe gpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(tap2apb_pclk_sync_rst_n),                                              // i:1
  .src_activity(glkp_activity),                                                 // i:1
  .src_strb(glkp_strb),                                                         // i:1
  .src_sop(glkp_sop),                                                           // i:1
  .src_eop(glkp_eop),                                                           // i:1
  .src_flitdata(glkp_flitdata),                                                 // i:36
  .src_ret_activity(glkp_ret_activity),                                         // o:1
  .src_ret_strb(glkp_ret_strb),                                                 // o:1
  .src_ret_cnt(glkp_ret_cnt),                                                   // o:1
  .dst_activity(glk_activity),                                                  // o:1
  .dst_strb(glk_strb),                                                          // o:1
  .dst_sop(glk_sop),                                                            // o:1
  .dst_eop(glk_eop),                                                            // o:1
  .dst_flitdata(glk_flitdata),                                                  // o:36
  .dst_ret_activity(glk_ret_activity),                                          // i:1
  .dst_ret_strb(glk_ret_strb),                                                  // i:1
  .dst_ret_cnt(glk_ret_cnt)                                                     // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_l2g_f0_lpipe lpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(llk_activity),                                                  // i:1
  .src_req(llk_req),                                                            // i:1
  .src_sop(llk_sop),                                                            // i:1
  .src_eop(llk_eop),                                                            // i:1
  .src_flitdata(llk_flitdata),                                                  // i:36
  .src_ready(llk_ready),                                                        // o:1
  .dst_activity(llkp_activity),                                                 // o:1
  .dst_req(llkp_req),                                                           // o:1
  .dst_sop(llkp_sop),                                                           // o:1
  .dst_eop(llkp_eop),                                                           // o:1
  .dst_flitdata(llkp_flitdata),                                                 // o:36
  .dst_ready(llkp_ready)                                                        // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_ls_l2g_f0_rstS rstS (
  .clk(tap2apb_pclk),                                                           // i:1
  .rawReset(tap2apb_pclk_sync_rst_n),                                           // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ========================================================
// Output Pipe
// ========================================================
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign glkp_activity = llkp_activity;
assign credclkEn = llkp_activity | glkp_ret_activity;
usb4_tc_noc_link0_ls_l2g_f0_creditcg creditcg (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(credclkEn),                                                            // i:1
  .clkOut(credclk),                                                             // o:1
  .isActive(credclkAct)                                                         // o:1
);
assign glkp_strb = llkp_req && llkp_ready;
assign glkp_flitdata = glkp_strb ? llkp_flitdata : 36'b0;
assign glkp_sop = glkp_strb ? llkp_sop      : 1'b0;
assign glkp_eop = glkp_strb ? llkp_eop      : 1'b0;
// Credit Tracking Logic
always_ff @(posedge credclk, negedge frst_n)
begin
  if (!frst_n)
    ccnt <= #1ps 12'd8;
  else if (ccnt_en)
    ccnt <= #1ps ccnt_nxt;
end

always_comb
begin
  ccnt_nxt = ccnt;
  ccnt_en = 1'b0;
  if (glkp_strb &&  glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt;                                           // 1's cancel out
      ccnt_en = 1'b1;
    end
  // We are transferring a flit and did not receive back credit in this cycle
  else if (glkp_strb)
    begin
      ccnt_nxt = ccnt - 1'd1;
      ccnt_en = 1'b1;
    end
  // We are not transferring a flit but did receive back credit  in this cycle
  else if (glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt + 1'd1;
      ccnt_en = 1'b1;
    end
end

assign llkp_ready = |(ccnt);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f0_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f0_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_ls_l2g_f0_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f0_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f0_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f0_creditcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f1 (
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  // llk
  input  wire            llk_activity,                                          // Upcoming activity indicator
  input  wire            llk_req,                                               // Flit transfer request
  input  wire            llk_sop,                                               // Start of packet indicator
  input  wire            llk_eop,                                               // End of packet indicator
  input  wire     [59:0] llk_flitdata,                                          // Flit data
  output logic           llk_ready,                                             // Flit transfer ready
  // glk
  output logic           glk_activity,                                          // Upcoming activity indicator
  output logic           glk_strb,                                              // Flit transfer strobe
  output logic           glk_sop,                                               // Start of Packet Flit Indicator
  output logic           glk_eop,                                               // End of Packet Flit Indicator
  output logic    [59:0] glk_flitdata,                                          // Flit data
  input  wire            glk_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            glk_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] glk_ret_cnt                                            // Credit return credit count
);

logic           glkp_activity;                                                  // Upcomong activity indicator
logic           glkp_strb;                                                      // Request
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [59:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [59:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           credclk;
logic           credclkAct;
wire            credclkEn;
logic    [11:0] ccnt;
logic    [11:0] ccnt_nxt;
logic     [0:0] ccnt_en;
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// LLK Interface
// ============================================
// ============================================
// LK Interface
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_l2g_f1_gpipe gpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(tap2apb_pclk_sync_rst_n),                                              // i:1
  .src_activity(glkp_activity),                                                 // i:1
  .src_strb(glkp_strb),                                                         // i:1
  .src_sop(glkp_sop),                                                           // i:1
  .src_eop(glkp_eop),                                                           // i:1
  .src_flitdata(glkp_flitdata),                                                 // i:60
  .src_ret_activity(glkp_ret_activity),                                         // o:1
  .src_ret_strb(glkp_ret_strb),                                                 // o:1
  .src_ret_cnt(glkp_ret_cnt),                                                   // o:1
  .dst_activity(glk_activity),                                                  // o:1
  .dst_strb(glk_strb),                                                          // o:1
  .dst_sop(glk_sop),                                                            // o:1
  .dst_eop(glk_eop),                                                            // o:1
  .dst_flitdata(glk_flitdata),                                                  // o:60
  .dst_ret_activity(glk_ret_activity),                                          // i:1
  .dst_ret_strb(glk_ret_strb),                                                  // i:1
  .dst_ret_cnt(glk_ret_cnt)                                                     // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_l2g_f1_lpipe lpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(llk_activity),                                                  // i:1
  .src_req(llk_req),                                                            // i:1
  .src_sop(llk_sop),                                                            // i:1
  .src_eop(llk_eop),                                                            // i:1
  .src_flitdata(llk_flitdata),                                                  // i:60
  .src_ready(llk_ready),                                                        // o:1
  .dst_activity(llkp_activity),                                                 // o:1
  .dst_req(llkp_req),                                                           // o:1
  .dst_sop(llkp_sop),                                                           // o:1
  .dst_eop(llkp_eop),                                                           // o:1
  .dst_flitdata(llkp_flitdata),                                                 // o:60
  .dst_ready(llkp_ready)                                                        // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_ls_l2g_f1_rstS rstS (
  .clk(tap2apb_pclk),                                                           // i:1
  .rawReset(tap2apb_pclk_sync_rst_n),                                           // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ========================================================
// Output Pipe
// ========================================================
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign glkp_activity = llkp_activity;
assign credclkEn = llkp_activity | glkp_ret_activity;
usb4_tc_noc_link0_ls_l2g_f1_creditcg creditcg (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(credclkEn),                                                            // i:1
  .clkOut(credclk),                                                             // o:1
  .isActive(credclkAct)                                                         // o:1
);
assign glkp_strb = llkp_req && llkp_ready;
assign glkp_flitdata = glkp_strb ? llkp_flitdata : 60'b0;
assign glkp_sop = glkp_strb ? llkp_sop      : 1'b0;
assign glkp_eop = glkp_strb ? llkp_eop      : 1'b0;
// Credit Tracking Logic
always_ff @(posedge credclk, negedge frst_n)
begin
  if (!frst_n)
    ccnt <= #1ps 12'd8;
  else if (ccnt_en)
    ccnt <= #1ps ccnt_nxt;
end

always_comb
begin
  ccnt_nxt = ccnt;
  ccnt_en = 1'b0;
  if (glkp_strb &&  glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt;                                           // 1's cancel out
      ccnt_en = 1'b1;
    end
  // We are transferring a flit and did not receive back credit in this cycle
  else if (glkp_strb)
    begin
      ccnt_nxt = ccnt - 1'd1;
      ccnt_en = 1'b1;
    end
  // We are not transferring a flit but did receive back credit  in this cycle
  else if (glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt + 1'd1;
      ccnt_en = 1'b1;
    end
end

assign llkp_ready = |(ccnt);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f1_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f1_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_ls_l2g_f1_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f1_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f1_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_l2g_f1_creditcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0 (
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  // glk
  input  wire            glk_activity,                                          // Upcomong activity indicator
  input  wire            glk_strb,                                              // Request
  input  wire            glk_sop,                                               // Start of Packet Flit Indicator
  input  wire            glk_eop,                                               // End of Packet Flit Indicator
  input  wire     [33:0] glk_flitdata,                                          // Flit data
  output logic           glk_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           glk_ret_strb,                                          // Credit return strobe
  output logic     [0:0] glk_ret_cnt,                                           // Credit return credit count
  // llk
  output logic           llk_activity,                                          // Upcoming activity indicator
  output logic           llk_req,                                               // Flit transfer request
  output logic           llk_sop,                                               // Start of packet indicator
  output logic           llk_eop,                                               // End of packet indicator
  output logic    [33:0] llk_flitdata,                                          // Flit data
  input  wire            llk_ready                                              // Flit transfer ready
);

logic           glkp_activity;                                                  // Upcoming activity indicator
logic           glkp_strb;                                                      // Flit transfer strobe
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [33:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [33:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           w_eop;                                                          // Write side eop
logic           wreq;                                                           // Write side req
logic    [33:0] wdata;                                                          // Write data
logic           wrdy;                                                           // Write side ready
logic           widle;                                                          // Valid on wclk
logic           cred_req;                                                       // Credit req
logic     [2:0] cred_val;                                                       // Credits transferred (credits-1)
logic           r_eop;                                                          // Read side eop
logic           rreq;                                                           // Read side req
logic           rrdy;                                                           // Read ready
logic           rrdy_active;                                                    // Read ready activity
logic    [33:0] rdata;                                                          // Read data
logic           Lfrst_n;                                                        // Output reset for async llk domain flops
logic           Llrst_n;                                                        // Output reset for everything else in llk domain
logic           Gfrst_n;                                                        // Output reset for async glk domain flops
logic           Glrst_n;                                                        // Output reset for everything else in glk domain
logic           gclkActive;                                                     // Activity synched to GLK clock
logic           gclkg;                                                          // GLK gated clock
logic           fwd_activity;                                                   // Forward activity synced to LLK clock
logic           rev_activity;                                                   // Reverse activity synced to GLK clock
logic           lclkActive;                                                     // Activity synched to LLK clock
logic           lclkg;                                                          // LLK gated clock
logic           gclkActiveSync;
logic     [0:0] gActive;
logic           rd;
logic     [0:0] inpkt;
logic           glkNotEmpty;
logic     [3:0] pendCred;
logic     [3:0] pendCred_nxt;
logic     [0:0] pendCred_en;
logic     [3:0] pendCredM1;
logic     [3:0] localReturn;
logic     [3:0] localRetCnt;
logic           llkNotEmpty;                                                    // We don't need help keeping the LLK side awake
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Credit Bus
// ============================================
// ============================================
// OCT Mode Tie-offs
// ============================================
// ============================================
// Global Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Local Port (LLK manager)
// ============================================
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_g2l_r0_gpipe gpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .src_activity(glk_activity),                                                  // i:1
  .src_strb(glk_strb),                                                          // i:1
  .src_sop(glk_sop),                                                            // i:1
  .src_eop(glk_eop),                                                            // i:1
  .src_flitdata(glk_flitdata),                                                  // i:34
  .src_ret_activity(glk_ret_activity),                                          // o:1
  .src_ret_strb(glk_ret_strb),                                                  // o:1
  .src_ret_cnt(glk_ret_cnt),                                                    // o:1
  .dst_activity(glkp_activity),                                                 // o:1
  .dst_strb(glkp_strb),                                                         // o:1
  .dst_sop(glkp_sop),                                                           // o:1
  .dst_eop(glkp_eop),                                                           // o:1
  .dst_flitdata(glkp_flitdata),                                                 // o:34
  .dst_ret_activity(glkp_ret_activity),                                         // i:1
  .dst_ret_strb(glkp_ret_strb),                                                 // i:1
  .dst_ret_cnt(glkp_ret_cnt)                                                    // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_g2l_r0_lpipe lpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .src_activity(llkp_activity),                                                 // i:1
  .src_req(llkp_req),                                                           // i:1
  .src_sop(llkp_sop),                                                           // i:1
  .src_eop(llkp_eop),                                                           // i:1
  .src_flitdata(llkp_flitdata),                                                 // i:34
  .src_ready(llkp_ready),                                                       // o:1
  .dst_activity(llk_activity),                                                  // o:1
  .dst_req(llk_req),                                                            // o:1
  .dst_sop(llk_sop),                                                            // o:1
  .dst_eop(llk_eop),                                                            // o:1
  .dst_flitdata(llk_flitdata),                                                  // o:34
  .dst_ready(llk_ready)                                                         // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_ls_g2l_r0_rstLS rstLS (
  .clk(tap2apb_pclk),                                                           // i:1
  .rawReset(tap2apb_pclk_sync_rst_n),                                           // i:1
  .flopReset(Lfrst_n),                                                          // o:1
  .logicReset(Llrst_n)                                                          // o:1
);
// If we have separate clocks, then we'll have separate sync'd resets,
// even if we only have a single reset coming into this module
usb4_tc_noc_link0_ls_g2l_r0_rstGS rstGS (
  .clk(noc_clk),                                                                // i:1
  .rawReset(noc_clk_sync_rst_n),                                                // i:1
  .flopReset(Gfrst_n),                                                          // o:1
  .logicReset(Glrst_n)                                                          // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_ls_g2l_r0_gclkcg gclkcg (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Gfrst_n),                                                              // i:1
  .enbIn(gclkActive),                                                           // i:1
  .clkOut(gclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Write side activity excludes read side
assign gclkActive = glkp_activity || glkNotEmpty || rev_activity;
// Async case: Flop the GLK side activity and synch it to the LLK side
always_ff @(posedge noc_clk, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    gActive <= #1ps 1'd0;
  else
    gActive <= #1ps gclkActive;
end

usb4_tc_noc_link0_ls_g2l_r0_activeSync activeSync (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .d(gActive),                                                                  // i:1
  .q(gclkActiveSync)                                                            // o:1
);
assign lclkActive = gclkActiveSync || llkNotEmpty;
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_ls_g2l_r0_lclkcg lclkcg (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .enbIn(lclkActive),                                                           // i:1
  .clkOut(lclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Send out our activity to our peers
assign glkp_ret_activity = rev_activity;
assign llkp_activity = fwd_activity;
// SOP generation
assign rd = llkp_req && llkp_ready;
always_ff @(posedge lclkg, negedge Lfrst_n)
begin
  if (!Lfrst_n)
    inpkt <= #1ps 1'd0;
  else if (rd)
    inpkt <= #1ps !llkp_eop;
end

assign llkp_sop = llkp_req && !inpkt;
usb4_tc_noc_link0_ls_g2l_r0_fifo fifo (
  .wclk(gclkg),                                                                 // i:1
  .w_rst_n(Gfrst_n),                                                            // i:1
  .rclk(lclkg),                                                                 // i:1
  .r_rst_n(Lfrst_n),                                                            // i:1
  .rclkSync(tap2apb_pclk),                                                      // i:1
  .w_eop(w_eop),                                                                // i:1
  .wreq(wreq),                                                                  // i:1
  .wdata(wdata),                                                                // i:34
  .wrdy(wrdy),                                                                  // o:1
  .widle(widle),                                                                // o:1
  .cred_req(cred_req),                                                          // o:1
  .cred_val(cred_val),                                                          // o:3
  .r_eop(r_eop),                                                                // o:1
  .rreq(rreq),                                                                  // i:1
  .rrdy(rrdy),                                                                  // o:1
  .rrdy_active(rrdy_active),                                                    // o:1
  .rdata(rdata)                                                                 // o:34
);
// GLK (Write) Side Logic
assign glkNotEmpty = !widle;
assign wreq = glkp_strb;
assign w_eop = glkp_eop;
assign wdata = glkp_flitdata;
always_ff @(posedge gclkg, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    pendCred <= #1ps 4'd0;
  else if (pendCred_en)
    pendCred <= #1ps pendCred_nxt;
end

always_comb
begin
  pendCred_nxt = pendCred;
  pendCred_en  = 1'b0;
  if( cred_req && glkp_ret_strb )
    begin
      pendCred_nxt = pendCred + cred_val - localRetCnt;                         // The 'd1 values cancel each other
      pendCred_en  = 1'b1;
    end
  else if( cred_req )
    begin
      pendCred_nxt = pendCred + cred_val + 4'd1;
      pendCred_en  = 1'b1;
    end
  else if( glkp_ret_strb )
    begin
      pendCred_nxt = pendCred - localRetCnt - 4'd1;
      pendCred_en  = 1'b1;
    end
end

assign rev_activity = |pendCred_nxt | glkp_ret_strb;
assign glkp_ret_strb = |pendCred;
assign pendCredM1 = pendCred - 4'd1;
assign localReturn = pendCred>4'd2 ? 4'd1 : pendCredM1;
assign localRetCnt = glkp_ret_strb ? localReturn : 4'd0;
assign glkp_ret_cnt = localRetCnt[0:0];
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// LLK (Read) Side Logic
assign fwd_activity = rrdy_active;
assign llkNotEmpty = 1'b0;                                                      // We don't need help keeping the LLK side awake
assign rreq = llkp_ready;
assign llkp_req = rrdy;
assign llkp_eop = r_eop;
assign llkp_flitdata = rdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_ls_g2l_r0_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_rstLS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_rstGS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_gclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_activeSync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [0:0] d,
  output wire      [0:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync (
  .xtout(q),                                                                    // (external)
  .xtin(d),                                                                     // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_lclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_fifo (
  input  wire            wclk,                                                  // Write side clock
  input  wire            w_rst_n,                                               // Write side reset
  input  wire            rclk,                                                  // Read side clock
  input  wire            r_rst_n,                                               // Read side reset
  input  wire            rclkSync,                                              // Read side clock (not gated)
  // write_side
  input  wire            w_eop,                                                 // Write side eop
  input  wire            wreq,                                                  // Write side req
  input  wire     [33:0] wdata,                                                 // Write data
  output logic           wrdy,                                                  // Write side ready
  output logic           widle,                                                 // Write side occupancy
  output logic           cred_req,                                              // Credit req
  output logic     [2:0] cred_val,                                              // Credits transferred (credits-1)
  // read_side
  output wire            r_eop,                                                 // Read side eop
  input  wire            rreq,                                                  // Read side req
  output wire            rrdy,                                                  // Read ready
  output wire            rrdy_active,                                           // Read ready activity
  output wire     [33:0] rdata                                                  // Read data
);

logic           put;
logic           get;
logic     [3:0] wp_ss_bin;
logic     [3:0] rp_ss_bin;
logic     [3:0] depth_wr;
logic     [3:0] depth_rd;
logic           full;                                                           // Valid on wclk
logic           empty;                                                          // Valid on rclk
logic     [2:0] waddr;
logic     [2:0] raddr;
logic           int_rrdy;
logic     [0:0] rrdy_enb;
logic     [3:0] rptrCred;
logic     [3:0] depth_credit;
logic     [2:0] creditm1;
logic     [3:0] wptr;
logic     [3:0] wptr_nxt;
logic     [0:0] wptr_en;
logic     [3:0] wptr_gray;
logic     [3:0] wptr_gray_nxt;
logic     [0:0] wptr_gray_en;
logic     [3:0] rptr;
logic     [3:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [3:0] rptr_gray;
logic     [3:0] rptr_gray_nxt;
logic     [0:0] rptr_gray_en;
logic     [3:0] rptr_gray_ss;
logic     [3:0] wptr_gray_ss;
logic    [34:0] sramRdata;
logic    [34:0] sramWdata;
// Ports
assign put = wreq && wrdy;
assign get = rreq && rrdy;
assign depth_wr = wptr - rp_ss_bin;
assign depth_rd = wp_ss_bin - rptr;
assign full = (depth_wr == 4'd8) ? 1'b1 : 1'b0;                                 // Valid on wclk
assign empty = (depth_rd == 4'd0) ? 1'b1 : 1'b0;                                // Valid on rclk
assign widle = (depth_wr == 4'd0) ? 1'b1 : 1'b0;                                // Valid on wclk
assign wrdy = !full;
assign r_eop = sramRdata[34];
assign rdata = sramRdata[33:0];
assign waddr = wptr[2:0];
assign raddr = rptr[2:0];
// Gray to binary
assign wp_ss_bin[0] = ^(wptr_gray_ss >> 2'd0);
assign rp_ss_bin[0] = ^(rptr_gray_ss >> 2'd0);
assign wp_ss_bin[1] = ^(wptr_gray_ss >> 2'd1);
assign rp_ss_bin[1] = ^(rptr_gray_ss >> 2'd1);
assign wp_ss_bin[2] = ^(wptr_gray_ss >> 2'd2);
assign rp_ss_bin[2] = ^(rptr_gray_ss >> 2'd2);
assign wp_ss_bin[3] = ^(wptr_gray_ss >> 2'd3);
assign rp_ss_bin[3] = ^(rptr_gray_ss >> 2'd3);
// Early rrdy logic
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rrdy_enb <= #1ps 1'd0;
  else
    rrdy_enb <= #1ps int_rrdy;
end

assign rrdy = int_rrdy && rrdy_enb;
assign rrdy_active = int_rrdy;
// Credit return
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    rptrCred <= #1ps 4'd0;
  else if (cred_req)
    rptrCred <= #1ps rp_ss_bin;
end

assign depth_credit = rp_ss_bin - rptrCred;
assign creditm1 = depth_credit[2:0] - 3'd1;
assign cred_val = creditm1;
assign cred_req = (|depth_credit);
// Write pointer / data
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr <= #1ps 4'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr_gray <= #1ps 4'd0;
  else if (wptr_gray_en)
    wptr_gray <= #1ps wptr_gray_nxt;
end

always_comb
begin
    wptr_nxt       = wptr;
    wptr_en        = 1'd0;
    wptr_gray_nxt  = wptr_gray;
    wptr_gray_en   = 1'd0;
    if (put)
        begin
            wptr_nxt        = wptr + 1'd1;
            wptr_en         = 1'd1;
            wptr_gray_nxt   = ((wptr + 1'd1)  >> 1) ^ (wptr + 1'd1);
            wptr_gray_en    = 1'd1;
        end
end

// Read Pointer
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr <= #1ps 4'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr_gray <= #1ps 4'd0;
  else if (rptr_gray_en)
    rptr_gray <= #1ps rptr_gray_nxt;
end

always_comb
begin
    rptr_nxt       = rptr;
    rptr_en        = 1'd0;
    rptr_gray_nxt  = rptr_gray;
    rptr_gray_en   = 1'd0;
    if (get)
        begin
            rptr_nxt =  rptr + 1'd1;
            rptr_en  = 1'd1;
            rptr_gray_nxt = ((rptr + 1'd1)  >> 1) ^ (rptr + 1'd1);
            rptr_gray_en  = 1'd1;
        end
end

// Synchronizers
usb4_tc_noc_link0_ls_g2l_r0_fifo_rsync rsync (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .d(rptr_gray),                                                                // i:4
  .q(rptr_gray_ss)                                                              // o:4
);
usb4_tc_noc_link0_ls_g2l_r0_fifo_wsync wsync (
  .clk(rclkSync),                                                               // i:1
  .rst_n(r_rst_n),                                                              // i:1
  .d(wptr_gray),                                                                // i:4
  .q(wptr_gray_ss)                                                              // o:4
);
// Data
assign sramWdata = {w_eop, wdata};
// Use a ansync read RAM
usb4_tc_noc_link0_ls_g2l_r0_fifo_fifoBuf fifoBuf (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .wen(put),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(sramWdata),                                                            // i:35
  .ren(rrdy),                                                                   // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(sramRdata)                                                             // o:35
);
// Optional holdback
assign int_rrdy = !empty;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_fifo_rsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_fifo_wsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r0_fifo_fifoBuf (
  input  wire            clk,
  input  wire            rst_n,
  // sramw
  input  wire            wen,
  input  wire      [2:0] waddr,
  input  wire     [34:0] wdata,
  // sramr
  input  wire            ren,
  input  wire      [2:0] raddr,
  output logic    [34:0] rdata
);

// tpRamCore Parameters
// Additional tpRam Parameters
usb4_tc_noc_tpRam_8_35_awn_raws usb4_tc_noc_tpRam_8_35_awn_raws (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .wen(wen),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(wdata),                                                                // i:35
  .ren(ren),                                                                    // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(rdata)                                                                 // o:35
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1 (
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  // glk
  input  wire            glk_activity,                                          // Upcomong activity indicator
  input  wire            glk_strb,                                              // Request
  input  wire            glk_sop,                                               // Start of Packet Flit Indicator
  input  wire            glk_eop,                                               // End of Packet Flit Indicator
  input  wire     [23:0] glk_flitdata,                                          // Flit data
  output logic           glk_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           glk_ret_strb,                                          // Credit return strobe
  output logic     [0:0] glk_ret_cnt,                                           // Credit return credit count
  // llk
  output logic           llk_activity,                                          // Upcoming activity indicator
  output logic           llk_req,                                               // Flit transfer request
  output logic           llk_sop,                                               // Start of packet indicator
  output logic           llk_eop,                                               // End of packet indicator
  output logic    [23:0] llk_flitdata,                                          // Flit data
  input  wire            llk_ready                                              // Flit transfer ready
);

logic           glkp_activity;                                                  // Upcoming activity indicator
logic           glkp_strb;                                                      // Flit transfer strobe
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [23:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [23:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           w_eop;                                                          // Write side eop
logic           wreq;                                                           // Write side req
logic    [23:0] wdata;                                                          // Write data
logic           wrdy;                                                           // Write side ready
logic           widle;                                                          // Valid on wclk
logic           cred_req;                                                       // Credit req
logic     [2:0] cred_val;                                                       // Credits transferred (credits-1)
logic           r_eop;                                                          // Read side eop
logic           rreq;                                                           // Read side req
logic           rrdy;                                                           // Read ready
logic           rrdy_active;                                                    // Read ready activity
logic    [23:0] rdata;                                                          // Read data
logic           Lfrst_n;                                                        // Output reset for async llk domain flops
logic           Llrst_n;                                                        // Output reset for everything else in llk domain
logic           Gfrst_n;                                                        // Output reset for async glk domain flops
logic           Glrst_n;                                                        // Output reset for everything else in glk domain
logic           gclkActive;                                                     // Activity synched to GLK clock
logic           gclkg;                                                          // GLK gated clock
logic           fwd_activity;                                                   // Forward activity synced to LLK clock
logic           rev_activity;                                                   // Reverse activity synced to GLK clock
logic           lclkActive;                                                     // Activity synched to LLK clock
logic           lclkg;                                                          // LLK gated clock
logic           gclkActiveSync;
logic     [0:0] gActive;
logic           rd;
logic     [0:0] inpkt;
logic           glkNotEmpty;
logic     [3:0] pendCred;
logic     [3:0] pendCred_nxt;
logic     [0:0] pendCred_en;
logic     [3:0] pendCredM1;
logic     [3:0] localReturn;
logic     [3:0] localRetCnt;
logic           llkNotEmpty;                                                    // We don't need help keeping the LLK side awake
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Credit Bus
// ============================================
// ============================================
// OCT Mode Tie-offs
// ============================================
// ============================================
// Global Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Local Port (LLK manager)
// ============================================
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_g2l_r1_gpipe gpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .src_activity(glk_activity),                                                  // i:1
  .src_strb(glk_strb),                                                          // i:1
  .src_sop(glk_sop),                                                            // i:1
  .src_eop(glk_eop),                                                            // i:1
  .src_flitdata(glk_flitdata),                                                  // i:24
  .src_ret_activity(glk_ret_activity),                                          // o:1
  .src_ret_strb(glk_ret_strb),                                                  // o:1
  .src_ret_cnt(glk_ret_cnt),                                                    // o:1
  .dst_activity(glkp_activity),                                                 // o:1
  .dst_strb(glkp_strb),                                                         // o:1
  .dst_sop(glkp_sop),                                                           // o:1
  .dst_eop(glkp_eop),                                                           // o:1
  .dst_flitdata(glkp_flitdata),                                                 // o:24
  .dst_ret_activity(glkp_ret_activity),                                         // i:1
  .dst_ret_strb(glkp_ret_strb),                                                 // i:1
  .dst_ret_cnt(glkp_ret_cnt)                                                    // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_ls_g2l_r1_lpipe lpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .src_activity(llkp_activity),                                                 // i:1
  .src_req(llkp_req),                                                           // i:1
  .src_sop(llkp_sop),                                                           // i:1
  .src_eop(llkp_eop),                                                           // i:1
  .src_flitdata(llkp_flitdata),                                                 // i:24
  .src_ready(llkp_ready),                                                       // o:1
  .dst_activity(llk_activity),                                                  // o:1
  .dst_req(llk_req),                                                            // o:1
  .dst_sop(llk_sop),                                                            // o:1
  .dst_eop(llk_eop),                                                            // o:1
  .dst_flitdata(llk_flitdata),                                                  // o:24
  .dst_ready(llk_ready)                                                         // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_ls_g2l_r1_rstLS rstLS (
  .clk(tap2apb_pclk),                                                           // i:1
  .rawReset(tap2apb_pclk_sync_rst_n),                                           // i:1
  .flopReset(Lfrst_n),                                                          // o:1
  .logicReset(Llrst_n)                                                          // o:1
);
// If we have separate clocks, then we'll have separate sync'd resets,
// even if we only have a single reset coming into this module
usb4_tc_noc_link0_ls_g2l_r1_rstGS rstGS (
  .clk(noc_clk),                                                                // i:1
  .rawReset(noc_clk_sync_rst_n),                                                // i:1
  .flopReset(Gfrst_n),                                                          // o:1
  .logicReset(Glrst_n)                                                          // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_ls_g2l_r1_gclkcg gclkcg (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Gfrst_n),                                                              // i:1
  .enbIn(gclkActive),                                                           // i:1
  .clkOut(gclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Write side activity excludes read side
assign gclkActive = glkp_activity || glkNotEmpty || rev_activity;
// Async case: Flop the GLK side activity and synch it to the LLK side
always_ff @(posedge noc_clk, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    gActive <= #1ps 1'd0;
  else
    gActive <= #1ps gclkActive;
end

usb4_tc_noc_link0_ls_g2l_r1_activeSync activeSync (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .d(gActive),                                                                  // i:1
  .q(gclkActiveSync)                                                            // o:1
);
assign lclkActive = gclkActiveSync || llkNotEmpty;
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_ls_g2l_r1_lclkcg lclkcg (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .enbIn(lclkActive),                                                           // i:1
  .clkOut(lclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Send out our activity to our peers
assign glkp_ret_activity = rev_activity;
assign llkp_activity = fwd_activity;
// SOP generation
assign rd = llkp_req && llkp_ready;
always_ff @(posedge lclkg, negedge Lfrst_n)
begin
  if (!Lfrst_n)
    inpkt <= #1ps 1'd0;
  else if (rd)
    inpkt <= #1ps !llkp_eop;
end

assign llkp_sop = llkp_req && !inpkt;
usb4_tc_noc_link0_ls_g2l_r1_fifo fifo (
  .wclk(gclkg),                                                                 // i:1
  .w_rst_n(Gfrst_n),                                                            // i:1
  .rclk(lclkg),                                                                 // i:1
  .r_rst_n(Lfrst_n),                                                            // i:1
  .rclkSync(tap2apb_pclk),                                                      // i:1
  .w_eop(w_eop),                                                                // i:1
  .wreq(wreq),                                                                  // i:1
  .wdata(wdata),                                                                // i:24
  .wrdy(wrdy),                                                                  // o:1
  .widle(widle),                                                                // o:1
  .cred_req(cred_req),                                                          // o:1
  .cred_val(cred_val),                                                          // o:3
  .r_eop(r_eop),                                                                // o:1
  .rreq(rreq),                                                                  // i:1
  .rrdy(rrdy),                                                                  // o:1
  .rrdy_active(rrdy_active),                                                    // o:1
  .rdata(rdata)                                                                 // o:24
);
// GLK (Write) Side Logic
assign glkNotEmpty = !widle;
assign wreq = glkp_strb;
assign w_eop = glkp_eop;
assign wdata = glkp_flitdata;
always_ff @(posedge gclkg, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    pendCred <= #1ps 4'd0;
  else if (pendCred_en)
    pendCred <= #1ps pendCred_nxt;
end

always_comb
begin
  pendCred_nxt = pendCred;
  pendCred_en  = 1'b0;
  if( cred_req && glkp_ret_strb )
    begin
      pendCred_nxt = pendCred + cred_val - localRetCnt;                         // The 'd1 values cancel each other
      pendCred_en  = 1'b1;
    end
  else if( cred_req )
    begin
      pendCred_nxt = pendCred + cred_val + 4'd1;
      pendCred_en  = 1'b1;
    end
  else if( glkp_ret_strb )
    begin
      pendCred_nxt = pendCred - localRetCnt - 4'd1;
      pendCred_en  = 1'b1;
    end
end

assign rev_activity = |pendCred_nxt | glkp_ret_strb;
assign glkp_ret_strb = |pendCred;
assign pendCredM1 = pendCred - 4'd1;
assign localReturn = pendCred>4'd2 ? 4'd1 : pendCredM1;
assign localRetCnt = glkp_ret_strb ? localReturn : 4'd0;
assign glkp_ret_cnt = localRetCnt[0:0];
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// LLK (Read) Side Logic
assign fwd_activity = rrdy_active;
assign llkNotEmpty = 1'b0;                                                      // We don't need help keeping the LLK side awake
assign rreq = llkp_ready;
assign llkp_req = rrdy;
assign llkp_eop = r_eop;
assign llkp_flitdata = rdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_ls_g2l_r1_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_rstLS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_rstGS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_gclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_activeSync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [0:0] d,
  output wire      [0:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync (
  .xtout(q),                                                                    // (external)
  .xtin(d),                                                                     // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_lclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_fifo (
  input  wire            wclk,                                                  // Write side clock
  input  wire            w_rst_n,                                               // Write side reset
  input  wire            rclk,                                                  // Read side clock
  input  wire            r_rst_n,                                               // Read side reset
  input  wire            rclkSync,                                              // Read side clock (not gated)
  // write_side
  input  wire            w_eop,                                                 // Write side eop
  input  wire            wreq,                                                  // Write side req
  input  wire     [23:0] wdata,                                                 // Write data
  output logic           wrdy,                                                  // Write side ready
  output logic           widle,                                                 // Write side occupancy
  output logic           cred_req,                                              // Credit req
  output logic     [2:0] cred_val,                                              // Credits transferred (credits-1)
  // read_side
  output wire            r_eop,                                                 // Read side eop
  input  wire            rreq,                                                  // Read side req
  output wire            rrdy,                                                  // Read ready
  output wire            rrdy_active,                                           // Read ready activity
  output wire     [23:0] rdata                                                  // Read data
);

logic           put;
logic           get;
logic     [3:0] wp_ss_bin;
logic     [3:0] rp_ss_bin;
logic     [3:0] depth_wr;
logic     [3:0] depth_rd;
logic           full;                                                           // Valid on wclk
logic           empty;                                                          // Valid on rclk
logic     [2:0] waddr;
logic     [2:0] raddr;
logic           int_rrdy;
logic     [0:0] rrdy_enb;
logic     [3:0] rptrCred;
logic     [3:0] depth_credit;
logic     [2:0] creditm1;
logic     [3:0] wptr;
logic     [3:0] wptr_nxt;
logic     [0:0] wptr_en;
logic     [3:0] wptr_gray;
logic     [3:0] wptr_gray_nxt;
logic     [0:0] wptr_gray_en;
logic     [3:0] rptr;
logic     [3:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [3:0] rptr_gray;
logic     [3:0] rptr_gray_nxt;
logic     [0:0] rptr_gray_en;
logic     [3:0] rptr_gray_ss;
logic     [3:0] wptr_gray_ss;
logic    [24:0] sramRdata;
logic    [24:0] sramWdata;
// Ports
assign put = wreq && wrdy;
assign get = rreq && rrdy;
assign depth_wr = wptr - rp_ss_bin;
assign depth_rd = wp_ss_bin - rptr;
assign full = (depth_wr == 4'd8) ? 1'b1 : 1'b0;                                 // Valid on wclk
assign empty = (depth_rd == 4'd0) ? 1'b1 : 1'b0;                                // Valid on rclk
assign widle = (depth_wr == 4'd0) ? 1'b1 : 1'b0;                                // Valid on wclk
assign wrdy = !full;
assign r_eop = sramRdata[24];
assign rdata = sramRdata[23:0];
assign waddr = wptr[2:0];
assign raddr = rptr[2:0];
// Gray to binary
assign wp_ss_bin[0] = ^(wptr_gray_ss >> 2'd0);
assign rp_ss_bin[0] = ^(rptr_gray_ss >> 2'd0);
assign wp_ss_bin[1] = ^(wptr_gray_ss >> 2'd1);
assign rp_ss_bin[1] = ^(rptr_gray_ss >> 2'd1);
assign wp_ss_bin[2] = ^(wptr_gray_ss >> 2'd2);
assign rp_ss_bin[2] = ^(rptr_gray_ss >> 2'd2);
assign wp_ss_bin[3] = ^(wptr_gray_ss >> 2'd3);
assign rp_ss_bin[3] = ^(rptr_gray_ss >> 2'd3);
// Early rrdy logic
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rrdy_enb <= #1ps 1'd0;
  else
    rrdy_enb <= #1ps int_rrdy;
end

assign rrdy = int_rrdy && rrdy_enb;
assign rrdy_active = int_rrdy;
// Credit return
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    rptrCred <= #1ps 4'd0;
  else if (cred_req)
    rptrCred <= #1ps rp_ss_bin;
end

assign depth_credit = rp_ss_bin - rptrCred;
assign creditm1 = depth_credit[2:0] - 3'd1;
assign cred_val = creditm1;
assign cred_req = (|depth_credit);
// Write pointer / data
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr <= #1ps 4'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr_gray <= #1ps 4'd0;
  else if (wptr_gray_en)
    wptr_gray <= #1ps wptr_gray_nxt;
end

always_comb
begin
    wptr_nxt       = wptr;
    wptr_en        = 1'd0;
    wptr_gray_nxt  = wptr_gray;
    wptr_gray_en   = 1'd0;
    if (put)
        begin
            wptr_nxt        = wptr + 1'd1;
            wptr_en         = 1'd1;
            wptr_gray_nxt   = ((wptr + 1'd1)  >> 1) ^ (wptr + 1'd1);
            wptr_gray_en    = 1'd1;
        end
end

// Read Pointer
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr <= #1ps 4'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr_gray <= #1ps 4'd0;
  else if (rptr_gray_en)
    rptr_gray <= #1ps rptr_gray_nxt;
end

always_comb
begin
    rptr_nxt       = rptr;
    rptr_en        = 1'd0;
    rptr_gray_nxt  = rptr_gray;
    rptr_gray_en   = 1'd0;
    if (get)
        begin
            rptr_nxt =  rptr + 1'd1;
            rptr_en  = 1'd1;
            rptr_gray_nxt = ((rptr + 1'd1)  >> 1) ^ (rptr + 1'd1);
            rptr_gray_en  = 1'd1;
        end
end

// Synchronizers
usb4_tc_noc_link0_ls_g2l_r1_fifo_rsync rsync (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .d(rptr_gray),                                                                // i:4
  .q(rptr_gray_ss)                                                              // o:4
);
usb4_tc_noc_link0_ls_g2l_r1_fifo_wsync wsync (
  .clk(rclkSync),                                                               // i:1
  .rst_n(r_rst_n),                                                              // i:1
  .d(wptr_gray),                                                                // i:4
  .q(wptr_gray_ss)                                                              // o:4
);
// Data
assign sramWdata = {w_eop, wdata};
// Use a ansync read RAM
usb4_tc_noc_link0_ls_g2l_r1_fifo_fifoBuf fifoBuf (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .wen(put),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(sramWdata),                                                            // i:25
  .ren(rrdy),                                                                   // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(sramRdata)                                                             // o:25
);
// Optional holdback
assign int_rrdy = !empty;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_fifo_rsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_fifo_wsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_ls_g2l_r1_fifo_fifoBuf (
  input  wire            clk,
  input  wire            rst_n,
  // sramw
  input  wire            wen,
  input  wire      [2:0] waddr,
  input  wire     [24:0] wdata,
  // sramr
  input  wire            ren,
  input  wire      [2:0] raddr,
  output logic    [24:0] rdata
);

// tpRamCore Parameters
// Additional tpRam Parameters
usb4_tc_noc_tpRam_8_25_awn_raws usb4_tc_noc_tpRam_8_25_awn_raws (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .wen(wen),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(wdata),                                                                // i:25
  .ren(ren),                                                                    // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(rdata)                                                                 // o:25
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt (
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  // glk_f0
  input  wire            glk_f0_activity,                                       // Upcomong activity indicator
  input  wire            glk_f0_strb,                                           // Request
  input  wire            glk_f0_sop,                                            // Start of Packet Flit Indicator
  input  wire            glk_f0_eop,                                            // End of Packet Flit Indicator
  input  wire     [35:0] glk_f0_flitdata,                                       // Flit data
  output logic           glk_f0_ret_activity,                                   // Upcoming credit return activity indicator
  output logic           glk_f0_ret_strb,                                       // Credit return strobe
  output logic     [0:0] glk_f0_ret_cnt,                                        // Credit return credit count
  // glk_f1
  input  wire            glk_f1_activity,                                       // Upcomong activity indicator
  input  wire            glk_f1_strb,                                           // Request
  input  wire            glk_f1_sop,                                            // Start of Packet Flit Indicator
  input  wire            glk_f1_eop,                                            // End of Packet Flit Indicator
  input  wire     [59:0] glk_f1_flitdata,                                       // Flit data
  output logic           glk_f1_ret_activity,                                   // Upcoming credit return activity indicator
  output logic           glk_f1_ret_strb,                                       // Credit return strobe
  output logic     [0:0] glk_f1_ret_cnt,                                        // Credit return credit count
  // glk_r0
  output logic           glk_r0_activity,                                       // Upcoming activity indicator
  output logic           glk_r0_strb,                                           // Flit transfer strobe
  output logic           glk_r0_sop,                                            // Start of Packet Flit Indicator
  output logic           glk_r0_eop,                                            // End of Packet Flit Indicator
  output logic    [33:0] glk_r0_flitdata,                                       // Flit data
  input  wire            glk_r0_ret_activity,                                   // Upcoming credit return activity indicator
  input  wire            glk_r0_ret_strb,                                       // Credit return strobe
  input  wire      [0:0] glk_r0_ret_cnt,                                        // Credit return credit count
  // glk_r1
  output logic           glk_r1_activity,                                       // Upcoming activity indicator
  output logic           glk_r1_strb,                                           // Flit transfer strobe
  output logic           glk_r1_sop,                                            // Start of Packet Flit Indicator
  output logic           glk_r1_eop,                                            // End of Packet Flit Indicator
  output logic    [23:0] glk_r1_flitdata,                                       // Flit data
  input  wire            glk_r1_ret_activity,                                   // Upcoming credit return activity indicator
  input  wire            glk_r1_ret_strb,                                       // Credit return strobe
  input  wire      [0:0] glk_r1_ret_cnt,                                        // Credit return credit count
  // llk_f0
  output logic           llk_f0_activity,                                       // Upcoming activity indicator
  output logic           llk_f0_req,                                            // Flit transfer request
  output logic           llk_f0_sop,                                            // Start of packet indicator
  output logic           llk_f0_eop,                                            // End of packet indicator
  output logic    [35:0] llk_f0_flitdata,                                       // Flit data
  input  wire            llk_f0_ready,                                          // Flit transfer ready
  // llk_f1
  output logic           llk_f1_activity,                                       // Upcoming activity indicator
  output logic           llk_f1_req,                                            // Flit transfer request
  output logic           llk_f1_sop,                                            // Start of packet indicator
  output logic           llk_f1_eop,                                            // End of packet indicator
  output logic    [59:0] llk_f1_flitdata,                                       // Flit data
  input  wire            llk_f1_ready,                                          // Flit transfer ready
  // llk_r0
  input  wire            llk_r0_activity,                                       // Upcoming activity indicator
  input  wire            llk_r0_req,                                            // Flit transfer request
  input  wire            llk_r0_sop,                                            // Start of packet indicator
  input  wire            llk_r0_eop,                                            // End of packet indicator
  input  wire     [33:0] llk_r0_flitdata,                                       // Flit data
  output logic           llk_r0_ready,                                          // Flit transfer ready
  // llk_r1
  input  wire            llk_r1_activity,                                       // Upcoming activity indicator
  input  wire            llk_r1_req,                                            // Flit transfer request
  input  wire            llk_r1_sop,                                            // Start of packet indicator
  input  wire            llk_r1_eop,                                            // End of packet indicator
  input  wire     [23:0] llk_r1_flitdata,                                       // Flit data
  output logic           llk_r1_ready                                           // Flit transfer ready
);

// =========================================================
// Clocks / Resets
// =========================================================
// Local clock / reset (may be only clock / reset)
// Global clock / reset
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// =========================================================
// Source Side LK Forward Channel Interfces (LK subordinate)
// =========================================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// =========================================================
// Source Side LLK Reverse Channel Interfaces (LK manager)
// =========================================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// =========================================================
// Dest Side LLK Forward Channel Interfaces (LLK manager)
// =========================================================
// =========================================================
// Dest Side LLK Reverse Channel Interfaces (LLK subordinate)
// =========================================================
// ===========================================
// NoC G2L Bridge Instances
// ===========================================
usb4_tc_noc_link0_lt_g2l_f0 g2l_f0 (
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .glk_activity(glk_f0_activity),                                               // i:1
  .glk_strb(glk_f0_strb),                                                       // i:1
  .glk_sop(glk_f0_sop),                                                         // i:1
  .glk_eop(glk_f0_eop),                                                         // i:1
  .glk_flitdata(glk_f0_flitdata),                                               // i:36
  .glk_ret_activity(glk_f0_ret_activity),                                       // o:1
  .glk_ret_strb(glk_f0_ret_strb),                                               // o:1
  .glk_ret_cnt(glk_f0_ret_cnt),                                                 // o:1
  .llk_activity(llk_f0_activity),                                               // o:1
  .llk_req(llk_f0_req),                                                         // o:1
  .llk_sop(llk_f0_sop),                                                         // o:1
  .llk_eop(llk_f0_eop),                                                         // o:1
  .llk_flitdata(llk_f0_flitdata),                                               // o:36
  .llk_ready(llk_f0_ready)                                                      // i:1
);
usb4_tc_noc_link0_lt_g2l_f1 g2l_f1 (
  .tap2apb_pclk(tap2apb_pclk),                                                  // i:1
  .tap2apb_pclk_sync_rst_n(tap2apb_pclk_sync_rst_n),                            // i:1
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .glk_activity(glk_f1_activity),                                               // i:1
  .glk_strb(glk_f1_strb),                                                       // i:1
  .glk_sop(glk_f1_sop),                                                         // i:1
  .glk_eop(glk_f1_eop),                                                         // i:1
  .glk_flitdata(glk_f1_flitdata),                                               // i:60
  .glk_ret_activity(glk_f1_ret_activity),                                       // o:1
  .glk_ret_strb(glk_f1_ret_strb),                                               // o:1
  .glk_ret_cnt(glk_f1_ret_cnt),                                                 // o:1
  .llk_activity(llk_f1_activity),                                               // o:1
  .llk_req(llk_f1_req),                                                         // o:1
  .llk_sop(llk_f1_sop),                                                         // o:1
  .llk_eop(llk_f1_eop),                                                         // o:1
  .llk_flitdata(llk_f1_flitdata),                                               // o:60
  .llk_ready(llk_f1_ready)                                                      // i:1
);
// ===========================================
// NoC G2L Bridge Instances
// ===========================================
usb4_tc_noc_link0_lt_l2g_r0 l2g_r0 (
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .llk_activity(llk_r0_activity),                                               // i:1
  .llk_req(llk_r0_req),                                                         // i:1
  .llk_sop(llk_r0_sop),                                                         // i:1
  .llk_eop(llk_r0_eop),                                                         // i:1
  .llk_flitdata(llk_r0_flitdata),                                               // i:34
  .llk_ready(llk_r0_ready),                                                     // o:1
  .glk_activity(glk_r0_activity),                                               // o:1
  .glk_strb(glk_r0_strb),                                                       // o:1
  .glk_sop(glk_r0_sop),                                                         // o:1
  .glk_eop(glk_r0_eop),                                                         // o:1
  .glk_flitdata(glk_r0_flitdata),                                               // o:34
  .glk_ret_activity(glk_r0_ret_activity),                                       // i:1
  .glk_ret_strb(glk_r0_ret_strb),                                               // i:1
  .glk_ret_cnt(glk_r0_ret_cnt)                                                  // i:1
);
usb4_tc_noc_link0_lt_l2g_r1 l2g_r1 (
  .noc_clk(noc_clk),                                                            // i:1
  .noc_clk_sync_rst_n(noc_clk_sync_rst_n),                                      // i:1
  .llk_activity(llk_r1_activity),                                               // i:1
  .llk_req(llk_r1_req),                                                         // i:1
  .llk_sop(llk_r1_sop),                                                         // i:1
  .llk_eop(llk_r1_eop),                                                         // i:1
  .llk_flitdata(llk_r1_flitdata),                                               // i:24
  .llk_ready(llk_r1_ready),                                                     // o:1
  .glk_activity(glk_r1_activity),                                               // o:1
  .glk_strb(glk_r1_strb),                                                       // o:1
  .glk_sop(glk_r1_sop),                                                         // o:1
  .glk_eop(glk_r1_eop),                                                         // o:1
  .glk_flitdata(glk_r1_flitdata),                                               // o:24
  .glk_ret_activity(glk_r1_ret_activity),                                       // i:1
  .glk_ret_strb(glk_r1_ret_strb),                                               // i:1
  .glk_ret_cnt(glk_r1_ret_cnt)                                                  // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0 (
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  // glk
  input  wire            glk_activity,                                          // Upcomong activity indicator
  input  wire            glk_strb,                                              // Request
  input  wire            glk_sop,                                               // Start of Packet Flit Indicator
  input  wire            glk_eop,                                               // End of Packet Flit Indicator
  input  wire     [35:0] glk_flitdata,                                          // Flit data
  output logic           glk_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           glk_ret_strb,                                          // Credit return strobe
  output logic     [0:0] glk_ret_cnt,                                           // Credit return credit count
  // llk
  output logic           llk_activity,                                          // Upcoming activity indicator
  output logic           llk_req,                                               // Flit transfer request
  output logic           llk_sop,                                               // Start of packet indicator
  output logic           llk_eop,                                               // End of packet indicator
  output logic    [35:0] llk_flitdata,                                          // Flit data
  input  wire            llk_ready                                              // Flit transfer ready
);

logic           glkp_activity;                                                  // Upcoming activity indicator
logic           glkp_strb;                                                      // Flit transfer strobe
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [35:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [35:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           w_eop;                                                          // Write side eop
logic           wreq;                                                           // Write side req
logic    [35:0] wdata;                                                          // Write data
logic           wrdy;                                                           // Write side ready
logic           widle;                                                          // Valid on wclk
logic           cred_req;                                                       // Credit req
logic     [2:0] cred_val;                                                       // Credits transferred (credits-1)
logic           r_eop;                                                          // Read side eop
logic           rreq;                                                           // Read side req
logic           rrdy;                                                           // Read ready
logic           rrdy_active;                                                    // Read ready activity
logic    [35:0] rdata;                                                          // Read data
logic           Lfrst_n;                                                        // Output reset for async llk domain flops
logic           Llrst_n;                                                        // Output reset for everything else in llk domain
logic           Gfrst_n;                                                        // Output reset for async glk domain flops
logic           Glrst_n;                                                        // Output reset for everything else in glk domain
logic           gclkActive;                                                     // Activity synched to GLK clock
logic           gclkg;                                                          // GLK gated clock
logic           fwd_activity;                                                   // Forward activity synced to LLK clock
logic           rev_activity;                                                   // Reverse activity synced to GLK clock
logic           lclkActive;                                                     // Activity synched to LLK clock
logic           lclkg;                                                          // LLK gated clock
logic           gclkActiveSync;
logic     [0:0] gActive;
logic           rd;
logic     [0:0] inpkt;
logic           glkNotEmpty;
logic     [3:0] pendCred;
logic     [3:0] pendCred_nxt;
logic     [0:0] pendCred_en;
logic     [3:0] pendCredM1;
logic     [3:0] localReturn;
logic     [3:0] localRetCnt;
logic           llkNotEmpty;                                                    // We don't need help keeping the LLK side awake
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Credit Bus
// ============================================
// ============================================
// OCT Mode Tie-offs
// ============================================
// ============================================
// Global Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Local Port (LLK manager)
// ============================================
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_g2l_f0_gpipe gpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(tap2apb_pclk_sync_rst_n),                                              // i:1
  .src_activity(glk_activity),                                                  // i:1
  .src_strb(glk_strb),                                                          // i:1
  .src_sop(glk_sop),                                                            // i:1
  .src_eop(glk_eop),                                                            // i:1
  .src_flitdata(glk_flitdata),                                                  // i:36
  .src_ret_activity(glk_ret_activity),                                          // o:1
  .src_ret_strb(glk_ret_strb),                                                  // o:1
  .src_ret_cnt(glk_ret_cnt),                                                    // o:1
  .dst_activity(glkp_activity),                                                 // o:1
  .dst_strb(glkp_strb),                                                         // o:1
  .dst_sop(glkp_sop),                                                           // o:1
  .dst_eop(glkp_eop),                                                           // o:1
  .dst_flitdata(glkp_flitdata),                                                 // o:36
  .dst_ret_activity(glkp_ret_activity),                                         // i:1
  .dst_ret_strb(glkp_ret_strb),                                                 // i:1
  .dst_ret_cnt(glkp_ret_cnt)                                                    // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_g2l_f0_lpipe lpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .src_activity(llkp_activity),                                                 // i:1
  .src_req(llkp_req),                                                           // i:1
  .src_sop(llkp_sop),                                                           // i:1
  .src_eop(llkp_eop),                                                           // i:1
  .src_flitdata(llkp_flitdata),                                                 // i:36
  .src_ready(llkp_ready),                                                       // o:1
  .dst_activity(llk_activity),                                                  // o:1
  .dst_req(llk_req),                                                            // o:1
  .dst_sop(llk_sop),                                                            // o:1
  .dst_eop(llk_eop),                                                            // o:1
  .dst_flitdata(llk_flitdata),                                                  // o:36
  .dst_ready(llk_ready)                                                         // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_lt_g2l_f0_rstLS rstLS (
  .clk(noc_clk),                                                                // i:1
  .rawReset(noc_clk_sync_rst_n),                                                // i:1
  .flopReset(Lfrst_n),                                                          // o:1
  .logicReset(Llrst_n)                                                          // o:1
);
// If we have separate clocks, then we'll have separate sync'd resets,
// even if we only have a single reset coming into this module
usb4_tc_noc_link0_lt_g2l_f0_rstGS rstGS (
  .clk(tap2apb_pclk),                                                           // i:1
  .rawReset(tap2apb_pclk_sync_rst_n),                                           // i:1
  .flopReset(Gfrst_n),                                                          // o:1
  .logicReset(Glrst_n)                                                          // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_lt_g2l_f0_gclkcg gclkcg (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Gfrst_n),                                                              // i:1
  .enbIn(gclkActive),                                                           // i:1
  .clkOut(gclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Write side activity excludes read side
assign gclkActive = glkp_activity || glkNotEmpty || rev_activity;
// Async case: Flop the GLK side activity and synch it to the LLK side
always_ff @(posedge tap2apb_pclk, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    gActive <= #1ps 1'd0;
  else
    gActive <= #1ps gclkActive;
end

usb4_tc_noc_link0_lt_g2l_f0_activeSync activeSync (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .d(gActive),                                                                  // i:1
  .q(gclkActiveSync)                                                            // o:1
);
assign lclkActive = gclkActiveSync || llkNotEmpty;
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_lt_g2l_f0_lclkcg lclkcg (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .enbIn(lclkActive),                                                           // i:1
  .clkOut(lclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Send out our activity to our peers
assign glkp_ret_activity = rev_activity;
assign llkp_activity = fwd_activity;
// SOP generation
assign rd = llkp_req && llkp_ready;
always_ff @(posedge lclkg, negedge Lfrst_n)
begin
  if (!Lfrst_n)
    inpkt <= #1ps 1'd0;
  else if (rd)
    inpkt <= #1ps !llkp_eop;
end

assign llkp_sop = llkp_req && !inpkt;
usb4_tc_noc_link0_lt_g2l_f0_fifo fifo (
  .wclk(gclkg),                                                                 // i:1
  .w_rst_n(Gfrst_n),                                                            // i:1
  .rclk(lclkg),                                                                 // i:1
  .r_rst_n(Lfrst_n),                                                            // i:1
  .rclkSync(noc_clk),                                                           // i:1
  .w_eop(w_eop),                                                                // i:1
  .wreq(wreq),                                                                  // i:1
  .wdata(wdata),                                                                // i:36
  .wrdy(wrdy),                                                                  // o:1
  .widle(widle),                                                                // o:1
  .cred_req(cred_req),                                                          // o:1
  .cred_val(cred_val),                                                          // o:3
  .r_eop(r_eop),                                                                // o:1
  .rreq(rreq),                                                                  // i:1
  .rrdy(rrdy),                                                                  // o:1
  .rrdy_active(rrdy_active),                                                    // o:1
  .rdata(rdata)                                                                 // o:36
);
// GLK (Write) Side Logic
assign glkNotEmpty = !widle;
assign wreq = glkp_strb;
assign w_eop = glkp_eop;
assign wdata = glkp_flitdata;
always_ff @(posedge gclkg, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    pendCred <= #1ps 4'd0;
  else if (pendCred_en)
    pendCred <= #1ps pendCred_nxt;
end

always_comb
begin
  pendCred_nxt = pendCred;
  pendCred_en  = 1'b0;
  if( cred_req && glkp_ret_strb )
    begin
      pendCred_nxt = pendCred + cred_val - localRetCnt;                         // The 'd1 values cancel each other
      pendCred_en  = 1'b1;
    end
  else if( cred_req )
    begin
      pendCred_nxt = pendCred + cred_val + 4'd1;
      pendCred_en  = 1'b1;
    end
  else if( glkp_ret_strb )
    begin
      pendCred_nxt = pendCred - localRetCnt - 4'd1;
      pendCred_en  = 1'b1;
    end
end

assign rev_activity = |pendCred_nxt | glkp_ret_strb;
assign glkp_ret_strb = |pendCred;
assign pendCredM1 = pendCred - 4'd1;
assign localReturn = pendCred>4'd2 ? 4'd1 : pendCredM1;
assign localRetCnt = glkp_ret_strb ? localReturn : 4'd0;
assign glkp_ret_cnt = localRetCnt[0:0];
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// LLK (Read) Side Logic
assign fwd_activity = rrdy_active;
assign llkNotEmpty = 1'b0;                                                      // We don't need help keeping the LLK side awake
assign rreq = llkp_ready;
assign llkp_req = rrdy;
assign llkp_eop = r_eop;
assign llkp_flitdata = rdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_lt_g2l_f0_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_rstLS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_rstGS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_gclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_activeSync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [0:0] d,
  output wire      [0:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync (
  .xtout(q),                                                                    // (external)
  .xtin(d),                                                                     // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_lclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_fifo (
  input  wire            wclk,                                                  // Write side clock
  input  wire            w_rst_n,                                               // Write side reset
  input  wire            rclk,                                                  // Read side clock
  input  wire            r_rst_n,                                               // Read side reset
  input  wire            rclkSync,                                              // Read side clock (not gated)
  // write_side
  input  wire            w_eop,                                                 // Write side eop
  input  wire            wreq,                                                  // Write side req
  input  wire     [35:0] wdata,                                                 // Write data
  output logic           wrdy,                                                  // Write side ready
  output logic           widle,                                                 // Write side occupancy
  output logic           cred_req,                                              // Credit req
  output logic     [2:0] cred_val,                                              // Credits transferred (credits-1)
  // read_side
  output wire            r_eop,                                                 // Read side eop
  input  wire            rreq,                                                  // Read side req
  output wire            rrdy,                                                  // Read ready
  output wire            rrdy_active,                                           // Read ready activity
  output wire     [35:0] rdata                                                  // Read data
);

logic           put;
logic           get;
logic     [3:0] wp_ss_bin;
logic     [3:0] rp_ss_bin;
logic     [3:0] depth_wr;
logic     [3:0] depth_rd;
logic           full;                                                           // Valid on wclk
logic           empty;                                                          // Valid on rclk
logic     [2:0] waddr;
logic     [2:0] raddr;
logic           int_rrdy;
logic     [0:0] rrdy_enb;
logic     [3:0] rptrCred;
logic     [3:0] depth_credit;
logic     [2:0] creditm1;
logic     [3:0] wptr;
logic     [3:0] wptr_nxt;
logic     [0:0] wptr_en;
logic     [3:0] wptr_gray;
logic     [3:0] wptr_gray_nxt;
logic     [0:0] wptr_gray_en;
logic     [3:0] rptr;
logic     [3:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [3:0] rptr_gray;
logic     [3:0] rptr_gray_nxt;
logic     [0:0] rptr_gray_en;
logic     [3:0] rptr_gray_ss;
logic     [3:0] wptr_gray_ss;
logic    [36:0] sramRdata;
logic    [36:0] sramWdata;
// Ports
assign put = wreq && wrdy;
assign get = rreq && rrdy;
assign depth_wr = wptr - rp_ss_bin;
assign depth_rd = wp_ss_bin - rptr;
assign full = (depth_wr == 4'd8) ? 1'b1 : 1'b0;                                 // Valid on wclk
assign empty = (depth_rd == 4'd0) ? 1'b1 : 1'b0;                                // Valid on rclk
assign widle = (depth_wr == 4'd0) ? 1'b1 : 1'b0;                                // Valid on wclk
assign wrdy = !full;
assign r_eop = sramRdata[36];
assign rdata = sramRdata[35:0];
assign waddr = wptr[2:0];
assign raddr = rptr[2:0];
// Gray to binary
assign wp_ss_bin[0] = ^(wptr_gray_ss >> 2'd0);
assign rp_ss_bin[0] = ^(rptr_gray_ss >> 2'd0);
assign wp_ss_bin[1] = ^(wptr_gray_ss >> 2'd1);
assign rp_ss_bin[1] = ^(rptr_gray_ss >> 2'd1);
assign wp_ss_bin[2] = ^(wptr_gray_ss >> 2'd2);
assign rp_ss_bin[2] = ^(rptr_gray_ss >> 2'd2);
assign wp_ss_bin[3] = ^(wptr_gray_ss >> 2'd3);
assign rp_ss_bin[3] = ^(rptr_gray_ss >> 2'd3);
// Early rrdy logic
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rrdy_enb <= #1ps 1'd0;
  else
    rrdy_enb <= #1ps int_rrdy;
end

assign rrdy = int_rrdy && rrdy_enb;
assign rrdy_active = int_rrdy;
// Credit return
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    rptrCred <= #1ps 4'd0;
  else if (cred_req)
    rptrCred <= #1ps rp_ss_bin;
end

assign depth_credit = rp_ss_bin - rptrCred;
assign creditm1 = depth_credit[2:0] - 3'd1;
assign cred_val = creditm1;
assign cred_req = (|depth_credit);
// Write pointer / data
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr <= #1ps 4'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr_gray <= #1ps 4'd0;
  else if (wptr_gray_en)
    wptr_gray <= #1ps wptr_gray_nxt;
end

always_comb
begin
    wptr_nxt       = wptr;
    wptr_en        = 1'd0;
    wptr_gray_nxt  = wptr_gray;
    wptr_gray_en   = 1'd0;
    if (put)
        begin
            wptr_nxt        = wptr + 1'd1;
            wptr_en         = 1'd1;
            wptr_gray_nxt   = ((wptr + 1'd1)  >> 1) ^ (wptr + 1'd1);
            wptr_gray_en    = 1'd1;
        end
end

// Read Pointer
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr <= #1ps 4'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr_gray <= #1ps 4'd0;
  else if (rptr_gray_en)
    rptr_gray <= #1ps rptr_gray_nxt;
end

always_comb
begin
    rptr_nxt       = rptr;
    rptr_en        = 1'd0;
    rptr_gray_nxt  = rptr_gray;
    rptr_gray_en   = 1'd0;
    if (get)
        begin
            rptr_nxt =  rptr + 1'd1;
            rptr_en  = 1'd1;
            rptr_gray_nxt = ((rptr + 1'd1)  >> 1) ^ (rptr + 1'd1);
            rptr_gray_en  = 1'd1;
        end
end

// Synchronizers
usb4_tc_noc_link0_lt_g2l_f0_fifo_rsync rsync (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .d(rptr_gray),                                                                // i:4
  .q(rptr_gray_ss)                                                              // o:4
);
usb4_tc_noc_link0_lt_g2l_f0_fifo_wsync wsync (
  .clk(rclkSync),                                                               // i:1
  .rst_n(r_rst_n),                                                              // i:1
  .d(wptr_gray),                                                                // i:4
  .q(wptr_gray_ss)                                                              // o:4
);
// Data
assign sramWdata = {w_eop, wdata};
// Use a ansync read RAM
usb4_tc_noc_link0_lt_g2l_f0_fifo_fifoBuf fifoBuf (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .wen(put),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(sramWdata),                                                            // i:37
  .ren(rrdy),                                                                   // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(sramRdata)                                                             // o:37
);
// Optional holdback
assign int_rrdy = !empty;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_fifo_rsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_fifo_wsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f0_fifo_fifoBuf (
  input  wire            clk,
  input  wire            rst_n,
  // sramw
  input  wire            wen,
  input  wire      [2:0] waddr,
  input  wire     [36:0] wdata,
  // sramr
  input  wire            ren,
  input  wire      [2:0] raddr,
  output logic    [36:0] rdata
);

// tpRamCore Parameters
// Additional tpRam Parameters
usb4_tc_noc_tpRam_8_37_awn_raws usb4_tc_noc_tpRam_8_37_awn_raws (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .wen(wen),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(wdata),                                                                // i:37
  .ren(ren),                                                                    // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(rdata)                                                                 // o:37
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1 (
  input  wire            tap2apb_pclk,
  input  wire            tap2apb_pclk_sync_rst_n,
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  // glk
  input  wire            glk_activity,                                          // Upcomong activity indicator
  input  wire            glk_strb,                                              // Request
  input  wire            glk_sop,                                               // Start of Packet Flit Indicator
  input  wire            glk_eop,                                               // End of Packet Flit Indicator
  input  wire     [59:0] glk_flitdata,                                          // Flit data
  output logic           glk_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           glk_ret_strb,                                          // Credit return strobe
  output logic     [0:0] glk_ret_cnt,                                           // Credit return credit count
  // llk
  output logic           llk_activity,                                          // Upcoming activity indicator
  output logic           llk_req,                                               // Flit transfer request
  output logic           llk_sop,                                               // Start of packet indicator
  output logic           llk_eop,                                               // End of packet indicator
  output logic    [59:0] llk_flitdata,                                          // Flit data
  input  wire            llk_ready                                              // Flit transfer ready
);

logic           glkp_activity;                                                  // Upcoming activity indicator
logic           glkp_strb;                                                      // Flit transfer strobe
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [59:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [59:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           w_eop;                                                          // Write side eop
logic           wreq;                                                           // Write side req
logic    [59:0] wdata;                                                          // Write data
logic           wrdy;                                                           // Write side ready
logic           widle;                                                          // Valid on wclk
logic           cred_req;                                                       // Credit req
logic     [2:0] cred_val;                                                       // Credits transferred (credits-1)
logic           r_eop;                                                          // Read side eop
logic           rreq;                                                           // Read side req
logic           rrdy;                                                           // Read ready
logic           rrdy_active;                                                    // Read ready activity
logic    [59:0] rdata;                                                          // Read data
logic           Lfrst_n;                                                        // Output reset for async llk domain flops
logic           Llrst_n;                                                        // Output reset for everything else in llk domain
logic           Gfrst_n;                                                        // Output reset for async glk domain flops
logic           Glrst_n;                                                        // Output reset for everything else in glk domain
logic           gclkActive;                                                     // Activity synched to GLK clock
logic           gclkg;                                                          // GLK gated clock
logic           fwd_activity;                                                   // Forward activity synced to LLK clock
logic           rev_activity;                                                   // Reverse activity synced to GLK clock
logic           lclkActive;                                                     // Activity synched to LLK clock
logic           lclkg;                                                          // LLK gated clock
logic           gclkActiveSync;
logic     [0:0] gActive;
logic           rd;
logic     [0:0] inpkt;
logic           glkNotEmpty;
logic     [3:0] pendCred;
logic     [3:0] pendCred_nxt;
logic     [0:0] pendCred_en;
logic     [3:0] pendCredM1;
logic     [3:0] localReturn;
logic     [3:0] localRetCnt;
logic           llkNotEmpty;                                                    // We don't need help keeping the LLK side awake
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Credit Bus
// ============================================
// ============================================
// OCT Mode Tie-offs
// ============================================
// ============================================
// Global Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Local Port (LLK manager)
// ============================================
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_g2l_f1_gpipe gpipe (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(tap2apb_pclk_sync_rst_n),                                              // i:1
  .src_activity(glk_activity),                                                  // i:1
  .src_strb(glk_strb),                                                          // i:1
  .src_sop(glk_sop),                                                            // i:1
  .src_eop(glk_eop),                                                            // i:1
  .src_flitdata(glk_flitdata),                                                  // i:60
  .src_ret_activity(glk_ret_activity),                                          // o:1
  .src_ret_strb(glk_ret_strb),                                                  // o:1
  .src_ret_cnt(glk_ret_cnt),                                                    // o:1
  .dst_activity(glkp_activity),                                                 // o:1
  .dst_strb(glkp_strb),                                                         // o:1
  .dst_sop(glkp_sop),                                                           // o:1
  .dst_eop(glkp_eop),                                                           // o:1
  .dst_flitdata(glkp_flitdata),                                                 // o:60
  .dst_ret_activity(glkp_ret_activity),                                         // i:1
  .dst_ret_strb(glkp_ret_strb),                                                 // i:1
  .dst_ret_cnt(glkp_ret_cnt)                                                    // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_g2l_f1_lpipe lpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .src_activity(llkp_activity),                                                 // i:1
  .src_req(llkp_req),                                                           // i:1
  .src_sop(llkp_sop),                                                           // i:1
  .src_eop(llkp_eop),                                                           // i:1
  .src_flitdata(llkp_flitdata),                                                 // i:60
  .src_ready(llkp_ready),                                                       // o:1
  .dst_activity(llk_activity),                                                  // o:1
  .dst_req(llk_req),                                                            // o:1
  .dst_sop(llk_sop),                                                            // o:1
  .dst_eop(llk_eop),                                                            // o:1
  .dst_flitdata(llk_flitdata),                                                  // o:60
  .dst_ready(llk_ready)                                                         // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_lt_g2l_f1_rstLS rstLS (
  .clk(noc_clk),                                                                // i:1
  .rawReset(noc_clk_sync_rst_n),                                                // i:1
  .flopReset(Lfrst_n),                                                          // o:1
  .logicReset(Llrst_n)                                                          // o:1
);
// If we have separate clocks, then we'll have separate sync'd resets,
// even if we only have a single reset coming into this module
usb4_tc_noc_link0_lt_g2l_f1_rstGS rstGS (
  .clk(tap2apb_pclk),                                                           // i:1
  .rawReset(tap2apb_pclk_sync_rst_n),                                           // i:1
  .flopReset(Gfrst_n),                                                          // o:1
  .logicReset(Glrst_n)                                                          // o:1
);
// ============================================
// Clock Gating Logic
// ============================================
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_lt_g2l_f1_gclkcg gclkcg (
  .clk(tap2apb_pclk),                                                           // i:1
  .rst_n(Gfrst_n),                                                              // i:1
  .enbIn(gclkActive),                                                           // i:1
  .clkOut(gclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Write side activity excludes read side
assign gclkActive = glkp_activity || glkNotEmpty || rev_activity;
// Async case: Flop the GLK side activity and synch it to the LLK side
always_ff @(posedge tap2apb_pclk, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    gActive <= #1ps 1'd0;
  else
    gActive <= #1ps gclkActive;
end

usb4_tc_noc_link0_lt_g2l_f1_activeSync activeSync (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .d(gActive),                                                                  // i:1
  .q(gclkActiveSync)                                                            // o:1
);
assign lclkActive = gclkActiveSync || llkNotEmpty;
// Use the activtity signal to gate the clock
usb4_tc_noc_link0_lt_g2l_f1_lclkcg lclkcg (
  .clk(noc_clk),                                                                // i:1
  .rst_n(Lfrst_n),                                                              // i:1
  .enbIn(lclkActive),                                                           // i:1
  .clkOut(lclkg),                                                               // o:1
  .isActive()                                                                   // o:1
);
// Send out our activity to our peers
assign glkp_ret_activity = rev_activity;
assign llkp_activity = fwd_activity;
// SOP generation
assign rd = llkp_req && llkp_ready;
always_ff @(posedge lclkg, negedge Lfrst_n)
begin
  if (!Lfrst_n)
    inpkt <= #1ps 1'd0;
  else if (rd)
    inpkt <= #1ps !llkp_eop;
end

assign llkp_sop = llkp_req && !inpkt;
usb4_tc_noc_link0_lt_g2l_f1_fifo fifo (
  .wclk(gclkg),                                                                 // i:1
  .w_rst_n(Gfrst_n),                                                            // i:1
  .rclk(lclkg),                                                                 // i:1
  .r_rst_n(Lfrst_n),                                                            // i:1
  .rclkSync(noc_clk),                                                           // i:1
  .w_eop(w_eop),                                                                // i:1
  .wreq(wreq),                                                                  // i:1
  .wdata(wdata),                                                                // i:60
  .wrdy(wrdy),                                                                  // o:1
  .widle(widle),                                                                // o:1
  .cred_req(cred_req),                                                          // o:1
  .cred_val(cred_val),                                                          // o:3
  .r_eop(r_eop),                                                                // o:1
  .rreq(rreq),                                                                  // i:1
  .rrdy(rrdy),                                                                  // o:1
  .rrdy_active(rrdy_active),                                                    // o:1
  .rdata(rdata)                                                                 // o:60
);
// GLK (Write) Side Logic
assign glkNotEmpty = !widle;
assign wreq = glkp_strb;
assign w_eop = glkp_eop;
assign wdata = glkp_flitdata;
always_ff @(posedge gclkg, negedge Gfrst_n)
begin
  if (!Gfrst_n)
    pendCred <= #1ps 4'd0;
  else if (pendCred_en)
    pendCred <= #1ps pendCred_nxt;
end

always_comb
begin
  pendCred_nxt = pendCred;
  pendCred_en  = 1'b0;
  if( cred_req && glkp_ret_strb )
    begin
      pendCred_nxt = pendCred + cred_val - localRetCnt;                         // The 'd1 values cancel each other
      pendCred_en  = 1'b1;
    end
  else if( cred_req )
    begin
      pendCred_nxt = pendCred + cred_val + 4'd1;
      pendCred_en  = 1'b1;
    end
  else if( glkp_ret_strb )
    begin
      pendCred_nxt = pendCred - localRetCnt - 4'd1;
      pendCred_en  = 1'b1;
    end
end

assign rev_activity = |pendCred_nxt | glkp_ret_strb;
assign glkp_ret_strb = |pendCred;
assign pendCredM1 = pendCred - 4'd1;
assign localReturn = pendCred>4'd2 ? 4'd1 : pendCredM1;
assign localRetCnt = glkp_ret_strb ? localReturn : 4'd0;
assign glkp_ret_cnt = localRetCnt[0:0];
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------------------------------------
// LLK (Read) Side Logic
assign fwd_activity = rrdy_active;
assign llkNotEmpty = 1'b0;                                                      // We don't need help keeping the LLK side awake
assign rreq = llkp_ready;
assign llkp_req = rrdy;
assign llkp_eop = r_eop;
assign llkp_flitdata = rdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_lt_g2l_f1_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_rstLS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_rstGS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_gclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_activeSync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [0:0] d,
  output wire      [0:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync (
  .xtout(q),                                                                    // (external)
  .xtin(d),                                                                     // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_lclkcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_fifo (
  input  wire            wclk,                                                  // Write side clock
  input  wire            w_rst_n,                                               // Write side reset
  input  wire            rclk,                                                  // Read side clock
  input  wire            r_rst_n,                                               // Read side reset
  input  wire            rclkSync,                                              // Read side clock (not gated)
  // write_side
  input  wire            w_eop,                                                 // Write side eop
  input  wire            wreq,                                                  // Write side req
  input  wire     [59:0] wdata,                                                 // Write data
  output logic           wrdy,                                                  // Write side ready
  output logic           widle,                                                 // Write side occupancy
  output logic           cred_req,                                              // Credit req
  output logic     [2:0] cred_val,                                              // Credits transferred (credits-1)
  // read_side
  output wire            r_eop,                                                 // Read side eop
  input  wire            rreq,                                                  // Read side req
  output wire            rrdy,                                                  // Read ready
  output wire            rrdy_active,                                           // Read ready activity
  output wire     [59:0] rdata                                                  // Read data
);

logic           put;
logic           get;
logic     [3:0] wp_ss_bin;
logic     [3:0] rp_ss_bin;
logic     [3:0] depth_wr;
logic     [3:0] depth_rd;
logic           full;                                                           // Valid on wclk
logic           empty;                                                          // Valid on rclk
logic     [2:0] waddr;
logic     [2:0] raddr;
logic           int_rrdy;
logic     [0:0] rrdy_enb;
logic     [3:0] rptrCred;
logic     [3:0] depth_credit;
logic     [2:0] creditm1;
logic     [3:0] wptr;
logic     [3:0] wptr_nxt;
logic     [0:0] wptr_en;
logic     [3:0] wptr_gray;
logic     [3:0] wptr_gray_nxt;
logic     [0:0] wptr_gray_en;
logic     [3:0] rptr;
logic     [3:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [3:0] rptr_gray;
logic     [3:0] rptr_gray_nxt;
logic     [0:0] rptr_gray_en;
logic     [3:0] rptr_gray_ss;
logic     [3:0] wptr_gray_ss;
logic    [60:0] sramRdata;
logic    [60:0] sramWdata;
// Ports
assign put = wreq && wrdy;
assign get = rreq && rrdy;
assign depth_wr = wptr - rp_ss_bin;
assign depth_rd = wp_ss_bin - rptr;
assign full = (depth_wr == 4'd8) ? 1'b1 : 1'b0;                                 // Valid on wclk
assign empty = (depth_rd == 4'd0) ? 1'b1 : 1'b0;                                // Valid on rclk
assign widle = (depth_wr == 4'd0) ? 1'b1 : 1'b0;                                // Valid on wclk
assign wrdy = !full;
assign r_eop = sramRdata[60];
assign rdata = sramRdata[59:0];
assign waddr = wptr[2:0];
assign raddr = rptr[2:0];
// Gray to binary
assign wp_ss_bin[0] = ^(wptr_gray_ss >> 2'd0);
assign rp_ss_bin[0] = ^(rptr_gray_ss >> 2'd0);
assign wp_ss_bin[1] = ^(wptr_gray_ss >> 2'd1);
assign rp_ss_bin[1] = ^(rptr_gray_ss >> 2'd1);
assign wp_ss_bin[2] = ^(wptr_gray_ss >> 2'd2);
assign rp_ss_bin[2] = ^(rptr_gray_ss >> 2'd2);
assign wp_ss_bin[3] = ^(wptr_gray_ss >> 2'd3);
assign rp_ss_bin[3] = ^(rptr_gray_ss >> 2'd3);
// Early rrdy logic
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rrdy_enb <= #1ps 1'd0;
  else
    rrdy_enb <= #1ps int_rrdy;
end

assign rrdy = int_rrdy && rrdy_enb;
assign rrdy_active = int_rrdy;
// Credit return
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    rptrCred <= #1ps 4'd0;
  else if (cred_req)
    rptrCred <= #1ps rp_ss_bin;
end

assign depth_credit = rp_ss_bin - rptrCred;
assign creditm1 = depth_credit[2:0] - 3'd1;
assign cred_val = creditm1;
assign cred_req = (|depth_credit);
// Write pointer / data
always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr <= #1ps 4'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_ff @(posedge wclk, negedge w_rst_n)
begin
  if (!w_rst_n)
    wptr_gray <= #1ps 4'd0;
  else if (wptr_gray_en)
    wptr_gray <= #1ps wptr_gray_nxt;
end

always_comb
begin
    wptr_nxt       = wptr;
    wptr_en        = 1'd0;
    wptr_gray_nxt  = wptr_gray;
    wptr_gray_en   = 1'd0;
    if (put)
        begin
            wptr_nxt        = wptr + 1'd1;
            wptr_en         = 1'd1;
            wptr_gray_nxt   = ((wptr + 1'd1)  >> 1) ^ (wptr + 1'd1);
            wptr_gray_en    = 1'd1;
        end
end

// Read Pointer
always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr <= #1ps 4'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_ff @(posedge rclk, negedge r_rst_n)
begin
  if (!r_rst_n)
    rptr_gray <= #1ps 4'd0;
  else if (rptr_gray_en)
    rptr_gray <= #1ps rptr_gray_nxt;
end

always_comb
begin
    rptr_nxt       = rptr;
    rptr_en        = 1'd0;
    rptr_gray_nxt  = rptr_gray;
    rptr_gray_en   = 1'd0;
    if (get)
        begin
            rptr_nxt =  rptr + 1'd1;
            rptr_en  = 1'd1;
            rptr_gray_nxt = ((rptr + 1'd1)  >> 1) ^ (rptr + 1'd1);
            rptr_gray_en  = 1'd1;
        end
end

// Synchronizers
usb4_tc_noc_link0_lt_g2l_f1_fifo_rsync rsync (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .d(rptr_gray),                                                                // i:4
  .q(rptr_gray_ss)                                                              // o:4
);
usb4_tc_noc_link0_lt_g2l_f1_fifo_wsync wsync (
  .clk(rclkSync),                                                               // i:1
  .rst_n(r_rst_n),                                                              // i:1
  .d(wptr_gray),                                                                // i:4
  .q(wptr_gray_ss)                                                              // o:4
);
// Data
assign sramWdata = {w_eop, wdata};
// Use a ansync read RAM
usb4_tc_noc_link0_lt_g2l_f1_fifo_fifoBuf fifoBuf (
  .clk(wclk),                                                                   // i:1
  .rst_n(w_rst_n),                                                              // i:1
  .wen(put),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(sramWdata),                                                            // i:61
  .ren(rrdy),                                                                   // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(sramRdata)                                                             // o:61
);
// Optional holdback
assign int_rrdy = !empty;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_fifo_rsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_fifo_wsync (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [3:0] d,
  output wire      [3:0] q
);

// Asynchronous Clear
// xtascsynch<N>( xtout, xtin, clrb, clk )
// Synchronous Clear
// xtscsynch<N>( xtout, xtin, clrb, clk )
// Non-Clearing
// xtsynch<N>( xtout, xtin, clk )
// Use asynch clear synchronizer
usb4_tc_noc_xtascsynch2 sync0 (
  .xtout(q[0]),                                                                 // (external)
  .xtin(d[0]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync1 (
  .xtout(q[1]),                                                                 // (external)
  .xtin(d[1]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync2 (
  .xtout(q[2]),                                                                 // (external)
  .xtin(d[2]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
usb4_tc_noc_xtascsynch2 sync3 (
  .xtout(q[3]),                                                                 // (external)
  .xtin(d[3]),                                                                  // (external)
  .clrb(rst_n),                                                                 // (external)
  .clk(clk)                                                                     // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_g2l_f1_fifo_fifoBuf (
  input  wire            clk,
  input  wire            rst_n,
  // sramw
  input  wire            wen,
  input  wire      [2:0] waddr,
  input  wire     [60:0] wdata,
  // sramr
  input  wire            ren,
  input  wire      [2:0] raddr,
  output logic    [60:0] rdata
);

// tpRamCore Parameters
// Additional tpRam Parameters
usb4_tc_noc_tpRam_8_61_awn_raws usb4_tc_noc_tpRam_8_61_awn_raws (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .wen(wen),                                                                    // i:1
  .waddr(waddr),                                                                // i:3
  .wdata(wdata),                                                                // i:61
  .ren(ren),                                                                    // i:1
  .raddr(raddr),                                                                // i:3
  .rdata(rdata)                                                                 // o:61
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r0 (
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  // llk
  input  wire            llk_activity,                                          // Upcoming activity indicator
  input  wire            llk_req,                                               // Flit transfer request
  input  wire            llk_sop,                                               // Start of packet indicator
  input  wire            llk_eop,                                               // End of packet indicator
  input  wire     [33:0] llk_flitdata,                                          // Flit data
  output logic           llk_ready,                                             // Flit transfer ready
  // glk
  output logic           glk_activity,                                          // Upcoming activity indicator
  output logic           glk_strb,                                              // Flit transfer strobe
  output logic           glk_sop,                                               // Start of Packet Flit Indicator
  output logic           glk_eop,                                               // End of Packet Flit Indicator
  output logic    [33:0] glk_flitdata,                                          // Flit data
  input  wire            glk_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            glk_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] glk_ret_cnt                                            // Credit return credit count
);

logic           glkp_activity;                                                  // Upcomong activity indicator
logic           glkp_strb;                                                      // Request
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [33:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [33:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           credclk;
logic           credclkAct;
wire            credclkEn;
logic    [11:0] ccnt;
logic    [11:0] ccnt_nxt;
logic     [0:0] ccnt_en;
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// LLK Interface
// ============================================
// ============================================
// LK Interface
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_l2g_r0_gpipe gpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .src_activity(glkp_activity),                                                 // i:1
  .src_strb(glkp_strb),                                                         // i:1
  .src_sop(glkp_sop),                                                           // i:1
  .src_eop(glkp_eop),                                                           // i:1
  .src_flitdata(glkp_flitdata),                                                 // i:34
  .src_ret_activity(glkp_ret_activity),                                         // o:1
  .src_ret_strb(glkp_ret_strb),                                                 // o:1
  .src_ret_cnt(glkp_ret_cnt),                                                   // o:1
  .dst_activity(glk_activity),                                                  // o:1
  .dst_strb(glk_strb),                                                          // o:1
  .dst_sop(glk_sop),                                                            // o:1
  .dst_eop(glk_eop),                                                            // o:1
  .dst_flitdata(glk_flitdata),                                                  // o:34
  .dst_ret_activity(glk_ret_activity),                                          // i:1
  .dst_ret_strb(glk_ret_strb),                                                  // i:1
  .dst_ret_cnt(glk_ret_cnt)                                                     // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_l2g_r0_lpipe lpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(llk_activity),                                                  // i:1
  .src_req(llk_req),                                                            // i:1
  .src_sop(llk_sop),                                                            // i:1
  .src_eop(llk_eop),                                                            // i:1
  .src_flitdata(llk_flitdata),                                                  // i:34
  .src_ready(llk_ready),                                                        // o:1
  .dst_activity(llkp_activity),                                                 // o:1
  .dst_req(llkp_req),                                                           // o:1
  .dst_sop(llkp_sop),                                                           // o:1
  .dst_eop(llkp_eop),                                                           // o:1
  .dst_flitdata(llkp_flitdata),                                                 // o:34
  .dst_ready(llkp_ready)                                                        // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_lt_l2g_r0_rstS rstS (
  .clk(noc_clk),                                                                // i:1
  .rawReset(noc_clk_sync_rst_n),                                                // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ========================================================
// Output Pipe
// ========================================================
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign glkp_activity = llkp_activity;
assign credclkEn = llkp_activity | glkp_ret_activity;
usb4_tc_noc_link0_lt_l2g_r0_creditcg creditcg (
  .clk(noc_clk),                                                                // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(credclkEn),                                                            // i:1
  .clkOut(credclk),                                                             // o:1
  .isActive(credclkAct)                                                         // o:1
);
assign glkp_strb = llkp_req && llkp_ready;
assign glkp_flitdata = glkp_strb ? llkp_flitdata : 34'b0;
assign glkp_sop = glkp_strb ? llkp_sop      : 1'b0;
assign glkp_eop = glkp_strb ? llkp_eop      : 1'b0;
// Credit Tracking Logic
always_ff @(posedge credclk, negedge frst_n)
begin
  if (!frst_n)
    ccnt <= #1ps 12'd8;
  else if (ccnt_en)
    ccnt <= #1ps ccnt_nxt;
end

always_comb
begin
  ccnt_nxt = ccnt;
  ccnt_en = 1'b0;
  if (glkp_strb &&  glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt;                                           // 1's cancel out
      ccnt_en = 1'b1;
    end
  // We are transferring a flit and did not receive back credit in this cycle
  else if (glkp_strb)
    begin
      ccnt_nxt = ccnt - 1'd1;
      ccnt_en = 1'b1;
    end
  // We are not transferring a flit but did receive back credit  in this cycle
  else if (glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt + 1'd1;
      ccnt_en = 1'b1;
    end
end

assign llkp_ready = |(ccnt);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r0_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r0_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_lt_l2g_r0_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r0_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r0_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r0_creditcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r1 (
  input  wire            noc_clk,
  input  wire            noc_clk_sync_rst_n,
  // llk
  input  wire            llk_activity,                                          // Upcoming activity indicator
  input  wire            llk_req,                                               // Flit transfer request
  input  wire            llk_sop,                                               // Start of packet indicator
  input  wire            llk_eop,                                               // End of packet indicator
  input  wire     [23:0] llk_flitdata,                                          // Flit data
  output logic           llk_ready,                                             // Flit transfer ready
  // glk
  output logic           glk_activity,                                          // Upcoming activity indicator
  output logic           glk_strb,                                              // Flit transfer strobe
  output logic           glk_sop,                                               // Start of Packet Flit Indicator
  output logic           glk_eop,                                               // End of Packet Flit Indicator
  output logic    [23:0] glk_flitdata,                                          // Flit data
  input  wire            glk_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            glk_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] glk_ret_cnt                                            // Credit return credit count
);

logic           glkp_activity;                                                  // Upcomong activity indicator
logic           glkp_strb;                                                      // Request
logic           glkp_sop;                                                       // Start of Packet Flit Indicator
logic           glkp_eop;                                                       // End of Packet Flit Indicator
logic    [23:0] glkp_flitdata;                                                  // Flit data
logic           glkp_ret_activity;                                              // Upcoming credit return activity indicator
logic           glkp_ret_strb;                                                  // Credit return strobe
logic     [0:0] glkp_ret_cnt;                                                   // Credit return credit count
logic           llkp_activity;                                                  // Upcoming activity indicator
logic           llkp_req;                                                       // Flit transfer request
logic           llkp_sop;                                                       // Start of packet indicator
logic           llkp_eop;                                                       // End of packet indicator
logic    [23:0] llkp_flitdata;                                                  // Flit data
logic           llkp_ready;                                                     // Flit transfer ready
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic           credclk;
logic           credclkAct;
wire            credclkEn;
logic    [11:0] ccnt;
logic    [11:0] ccnt_nxt;
logic     [0:0] ccnt_en;
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// LLK Interface
// ============================================
// ============================================
// LK Interface
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Global Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_l2g_r1_gpipe gpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(noc_clk_sync_rst_n),                                                   // i:1
  .src_activity(glkp_activity),                                                 // i:1
  .src_strb(glkp_strb),                                                         // i:1
  .src_sop(glkp_sop),                                                           // i:1
  .src_eop(glkp_eop),                                                           // i:1
  .src_flitdata(glkp_flitdata),                                                 // i:24
  .src_ret_activity(glkp_ret_activity),                                         // o:1
  .src_ret_strb(glkp_ret_strb),                                                 // o:1
  .src_ret_cnt(glkp_ret_cnt),                                                   // o:1
  .dst_activity(glk_activity),                                                  // o:1
  .dst_strb(glk_strb),                                                          // o:1
  .dst_sop(glk_sop),                                                            // o:1
  .dst_eop(glk_eop),                                                            // o:1
  .dst_flitdata(glk_flitdata),                                                  // o:24
  .dst_ret_activity(glk_ret_activity),                                          // i:1
  .dst_ret_strb(glk_ret_strb),                                                  // i:1
  .dst_ret_cnt(glk_ret_cnt)                                                     // i:1
);
// ============================================
// Local Link Interface Pipe Stage
// ============================================
usb4_tc_noc_link0_lt_l2g_r1_lpipe lpipe (
  .clk(noc_clk),                                                                // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(llk_activity),                                                  // i:1
  .src_req(llk_req),                                                            // i:1
  .src_sop(llk_sop),                                                            // i:1
  .src_eop(llk_eop),                                                            // i:1
  .src_flitdata(llk_flitdata),                                                  // i:24
  .src_ready(llk_ready),                                                        // o:1
  .dst_activity(llkp_activity),                                                 // o:1
  .dst_req(llkp_req),                                                           // o:1
  .dst_sop(llkp_sop),                                                           // o:1
  .dst_eop(llkp_eop),                                                           // o:1
  .dst_flitdata(llkp_flitdata),                                                 // o:24
  .dst_ready(llkp_ready)                                                        // i:1
);
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_link0_lt_l2g_r1_rstS rstS (
  .clk(noc_clk),                                                                // i:1
  .rawReset(noc_clk_sync_rst_n),                                                // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ========================================================
// Output Pipe
// ========================================================
// ============================================
// Clock Gating Logic
// ============================================
// APB state clock
assign glkp_activity = llkp_activity;
assign credclkEn = llkp_activity | glkp_ret_activity;
usb4_tc_noc_link0_lt_l2g_r1_creditcg creditcg (
  .clk(noc_clk),                                                                // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(credclkEn),                                                            // i:1
  .clkOut(credclk),                                                             // o:1
  .isActive(credclkAct)                                                         // o:1
);
assign glkp_strb = llkp_req && llkp_ready;
assign glkp_flitdata = glkp_strb ? llkp_flitdata : 24'b0;
assign glkp_sop = glkp_strb ? llkp_sop      : 1'b0;
assign glkp_eop = glkp_strb ? llkp_eop      : 1'b0;
// Credit Tracking Logic
always_ff @(posedge credclk, negedge frst_n)
begin
  if (!frst_n)
    ccnt <= #1ps 12'd8;
  else if (ccnt_en)
    ccnt <= #1ps ccnt_nxt;
end

always_comb
begin
  ccnt_nxt = ccnt;
  ccnt_en = 1'b0;
  if (glkp_strb &&  glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt;                                           // 1's cancel out
      ccnt_en = 1'b1;
    end
  // We are transferring a flit and did not receive back credit in this cycle
  else if (glkp_strb)
    begin
      ccnt_nxt = ccnt - 1'd1;
      ccnt_en = 1'b1;
    end
  // We are not transferring a flit but did receive back credit  in this cycle
  else if (glkp_ret_strb)
    begin
      ccnt_nxt = ccnt + glkp_ret_cnt + 1'd1;
      ccnt_en = 1'b1;
    end
end

assign llkp_ready = |(ccnt);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r1_gpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcomong activity indicator
  input  wire            src_strb,                                              // Request
  input  wire            src_sop,                                               // Start of Packet Flit Indicator
  input  wire            src_eop,                                               // End of Packet Flit Indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ret_activity,                                      // Upcoming credit return activity indicator
  output logic           src_ret_strb,                                          // Credit return strobe
  output logic     [0:0] src_ret_cnt,                                           // Credit return credit count
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_strb,                                              // Flit transfer strobe
  output logic           dst_sop,                                               // Start of Packet Flit Indicator
  output logic           dst_eop,                                               // End of Packet Flit Indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ret_activity,                                      // Upcoming credit return activity indicator
  input  wire            dst_ret_strb,                                          // Credit return strobe
  input  wire      [0:0] dst_ret_cnt                                            // Credit return credit count
);

// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LK subordinate)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ============================================
// Destination Port (LK manager)
// ============================================
// Manager view of pins
// Subordinate view of pins
// Monitor view of pins
// Bus view of pins (internal interface within module)
// ===========================================
// Outputs
// ===========================================
assign dst_activity = src_activity;
assign src_ret_activity = dst_ret_activity;
assign dst_strb = src_strb;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
assign src_ret_strb = dst_ret_strb;
assign src_ret_cnt = dst_ret_cnt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r1_lpipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_link0_lt_l2g_r1_lpipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r1_lpipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r1_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_link0_lt_l2g_r1_creditcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0 (
  input  wire            clk,
  input  wire            rst_n,
  // apb_mstr_f0
  input  wire            apb_mstr_f0_activity,                                  // Upcoming activity indicator
  input  wire            apb_mstr_f0_req,                                       // Flit transfer request
  input  wire            apb_mstr_f0_sop,                                       // Start of packet indicator
  input  wire            apb_mstr_f0_eop,                                       // End of packet indicator
  input  wire     [35:0] apb_mstr_f0_flitdata,                                  // Flit data
  output logic           apb_mstr_f0_ready,                                     // Flit transfer ready
  // apb_mstr_f1
  input  wire            apb_mstr_f1_activity,                                  // Upcoming activity indicator
  input  wire            apb_mstr_f1_req,                                       // Flit transfer request
  input  wire            apb_mstr_f1_sop,                                       // Start of packet indicator
  input  wire            apb_mstr_f1_eop,                                       // End of packet indicator
  input  wire     [59:0] apb_mstr_f1_flitdata,                                  // Flit data
  output logic           apb_mstr_f1_ready,                                     // Flit transfer ready
  // apb_mstr_r0
  output logic           apb_mstr_r0_activity,                                  // Upcoming activity indicator
  output logic           apb_mstr_r0_req,                                       // Flit transfer request
  output logic           apb_mstr_r0_sop,                                       // Start of packet indicator
  output logic           apb_mstr_r0_eop,                                       // End of packet indicator
  output logic    [33:0] apb_mstr_r0_flitdata,                                  // Flit data
  input  wire            apb_mstr_r0_ready,                                     // Flit transfer ready
  // apb_mstr_r1
  output logic           apb_mstr_r1_activity,                                  // Upcoming activity indicator
  output logic           apb_mstr_r1_req,                                       // Flit transfer request
  output logic           apb_mstr_r1_sop,                                       // Start of packet indicator
  output logic           apb_mstr_r1_eop,                                       // End of packet indicator
  output logic    [23:0] apb_mstr_r1_flitdata,                                  // Flit data
  input  wire            apb_mstr_r1_ready,                                     // Flit transfer ready
  // RTR_INI0_f0
  input  wire            RTR_INI0_f0_activity,                                  // Upcoming activity indicator
  input  wire            RTR_INI0_f0_req,                                       // Flit transfer request
  input  wire            RTR_INI0_f0_sop,                                       // Start of packet indicator
  input  wire            RTR_INI0_f0_eop,                                       // End of packet indicator
  input  wire     [35:0] RTR_INI0_f0_flitdata,                                  // Flit data
  output logic           RTR_INI0_f0_ready,                                     // Flit transfer ready
  // RTR_INI0_f1
  input  wire            RTR_INI0_f1_activity,                                  // Upcoming activity indicator
  input  wire            RTR_INI0_f1_req,                                       // Flit transfer request
  input  wire            RTR_INI0_f1_sop,                                       // Start of packet indicator
  input  wire            RTR_INI0_f1_eop,                                       // End of packet indicator
  input  wire     [59:0] RTR_INI0_f1_flitdata,                                  // Flit data
  output logic           RTR_INI0_f1_ready,                                     // Flit transfer ready
  // RTR_INI0_r0
  output logic           RTR_INI0_r0_activity,                                  // Upcoming activity indicator
  output logic           RTR_INI0_r0_req,                                       // Flit transfer request
  output logic           RTR_INI0_r0_sop,                                       // Start of packet indicator
  output logic           RTR_INI0_r0_eop,                                       // End of packet indicator
  output logic    [33:0] RTR_INI0_r0_flitdata,                                  // Flit data
  input  wire            RTR_INI0_r0_ready,                                     // Flit transfer ready
  // RTR_INI0_r1
  output logic           RTR_INI0_r1_activity,                                  // Upcoming activity indicator
  output logic           RTR_INI0_r1_req,                                       // Flit transfer request
  output logic           RTR_INI0_r1_sop,                                       // Start of packet indicator
  output logic           RTR_INI0_r1_eop,                                       // End of packet indicator
  output logic    [23:0] RTR_INI0_r1_flitdata,                                  // Flit data
  input  wire            RTR_INI0_r1_ready,                                     // Flit transfer ready
  // pam3_cmn_TEA_f0
  output logic           pam3_cmn_TEA_f0_activity,                              // Upcoming activity indicator
  output logic           pam3_cmn_TEA_f0_req,                                   // Flit transfer request
  output logic           pam3_cmn_TEA_f0_sop,                                   // Start of packet indicator
  output logic           pam3_cmn_TEA_f0_eop,                                   // End of packet indicator
  output logic    [35:0] pam3_cmn_TEA_f0_flitdata,                              // Flit data
  input  wire            pam3_cmn_TEA_f0_ready,                                 // Flit transfer ready
  // pam3_cmn_TEA_f1
  output logic           pam3_cmn_TEA_f1_activity,                              // Upcoming activity indicator
  output logic           pam3_cmn_TEA_f1_req,                                   // Flit transfer request
  output logic           pam3_cmn_TEA_f1_sop,                                   // Start of packet indicator
  output logic           pam3_cmn_TEA_f1_eop,                                   // End of packet indicator
  output logic    [59:0] pam3_cmn_TEA_f1_flitdata,                              // Flit data
  input  wire            pam3_cmn_TEA_f1_ready,                                 // Flit transfer ready
  // pam3_cmn_TEA_r0
  input  wire            pam3_cmn_TEA_r0_activity,                              // Upcoming activity indicator
  input  wire            pam3_cmn_TEA_r0_req,                                   // Flit transfer request
  input  wire            pam3_cmn_TEA_r0_sop,                                   // Start of packet indicator
  input  wire            pam3_cmn_TEA_r0_eop,                                   // End of packet indicator
  input  wire     [33:0] pam3_cmn_TEA_r0_flitdata,                              // Flit data
  output logic           pam3_cmn_TEA_r0_ready,                                 // Flit transfer ready
  // pam3_cmn_TEA_r1
  input  wire            pam3_cmn_TEA_r1_activity,                              // Upcoming activity indicator
  input  wire            pam3_cmn_TEA_r1_req,                                   // Flit transfer request
  input  wire            pam3_cmn_TEA_r1_sop,                                   // Start of packet indicator
  input  wire            pam3_cmn_TEA_r1_eop,                                   // End of packet indicator
  input  wire     [23:0] pam3_cmn_TEA_r1_flitdata,                              // Flit data
  output logic           pam3_cmn_TEA_r1_ready,                                 // Flit transfer ready
  // tc_reg_TEA_f0
  output logic           tc_reg_TEA_f0_activity,                                // Upcoming activity indicator
  output logic           tc_reg_TEA_f0_req,                                     // Flit transfer request
  output logic           tc_reg_TEA_f0_sop,                                     // Start of packet indicator
  output logic           tc_reg_TEA_f0_eop,                                     // End of packet indicator
  output logic    [35:0] tc_reg_TEA_f0_flitdata,                                // Flit data
  input  wire            tc_reg_TEA_f0_ready,                                   // Flit transfer ready
  // tc_reg_TEA_f1
  output logic           tc_reg_TEA_f1_activity,                                // Upcoming activity indicator
  output logic           tc_reg_TEA_f1_req,                                     // Flit transfer request
  output logic           tc_reg_TEA_f1_sop,                                     // Start of packet indicator
  output logic           tc_reg_TEA_f1_eop,                                     // End of packet indicator
  output logic    [59:0] tc_reg_TEA_f1_flitdata,                                // Flit data
  input  wire            tc_reg_TEA_f1_ready,                                   // Flit transfer ready
  // tc_reg_TEA_r0
  input  wire            tc_reg_TEA_r0_activity,                                // Upcoming activity indicator
  input  wire            tc_reg_TEA_r0_req,                                     // Flit transfer request
  input  wire            tc_reg_TEA_r0_sop,                                     // Start of packet indicator
  input  wire            tc_reg_TEA_r0_eop,                                     // End of packet indicator
  input  wire     [33:0] tc_reg_TEA_r0_flitdata,                                // Flit data
  output logic           tc_reg_TEA_r0_ready,                                   // Flit transfer ready
  // tc_reg_TEA_r1
  input  wire            tc_reg_TEA_r1_activity,                                // Upcoming activity indicator
  input  wire            tc_reg_TEA_r1_req,                                     // Flit transfer request
  input  wire            tc_reg_TEA_r1_sop,                                     // Start of packet indicator
  input  wire            tc_reg_TEA_r1_eop,                                     // End of packet indicator
  input  wire     [23:0] tc_reg_TEA_r1_flitdata,                                // Flit data
  output logic           tc_reg_TEA_r1_ready,                                   // Flit transfer ready
  // usb_sub_sys_TEA_f0
  output logic           usb_sub_sys_TEA_f0_activity,                           // Upcoming activity indicator
  output logic           usb_sub_sys_TEA_f0_req,                                // Flit transfer request
  output logic           usb_sub_sys_TEA_f0_sop,                                // Start of packet indicator
  output logic           usb_sub_sys_TEA_f0_eop,                                // End of packet indicator
  output logic    [35:0] usb_sub_sys_TEA_f0_flitdata,                           // Flit data
  input  wire            usb_sub_sys_TEA_f0_ready,                              // Flit transfer ready
  // usb_sub_sys_TEA_f1
  output logic           usb_sub_sys_TEA_f1_activity,                           // Upcoming activity indicator
  output logic           usb_sub_sys_TEA_f1_req,                                // Flit transfer request
  output logic           usb_sub_sys_TEA_f1_sop,                                // Start of packet indicator
  output logic           usb_sub_sys_TEA_f1_eop,                                // End of packet indicator
  output logic    [59:0] usb_sub_sys_TEA_f1_flitdata,                           // Flit data
  input  wire            usb_sub_sys_TEA_f1_ready,                              // Flit transfer ready
  // usb_sub_sys_TEA_r0
  input  wire            usb_sub_sys_TEA_r0_activity,                           // Upcoming activity indicator
  input  wire            usb_sub_sys_TEA_r0_req,                                // Flit transfer request
  input  wire            usb_sub_sys_TEA_r0_sop,                                // Start of packet indicator
  input  wire            usb_sub_sys_TEA_r0_eop,                                // End of packet indicator
  input  wire     [33:0] usb_sub_sys_TEA_r0_flitdata,                           // Flit data
  output logic           usb_sub_sys_TEA_r0_ready,                              // Flit transfer ready
  // usb_sub_sys_TEA_r1
  input  wire            usb_sub_sys_TEA_r1_activity,                           // Upcoming activity indicator
  input  wire            usb_sub_sys_TEA_r1_req,                                // Flit transfer request
  input  wire            usb_sub_sys_TEA_r1_sop,                                // Start of packet indicator
  input  wire            usb_sub_sys_TEA_r1_eop,                                // End of packet indicator
  input  wire     [23:0] usb_sub_sys_TEA_r1_flitdata,                           // Flit data
  output logic           usb_sub_sys_TEA_r1_ready,                              // Flit transfer ready
  // pam3_sub_sys_TEA_f0
  output logic           pam3_sub_sys_TEA_f0_activity,                          // Upcoming activity indicator
  output logic           pam3_sub_sys_TEA_f0_req,                               // Flit transfer request
  output logic           pam3_sub_sys_TEA_f0_sop,                               // Start of packet indicator
  output logic           pam3_sub_sys_TEA_f0_eop,                               // End of packet indicator
  output logic    [35:0] pam3_sub_sys_TEA_f0_flitdata,                          // Flit data
  input  wire            pam3_sub_sys_TEA_f0_ready,                             // Flit transfer ready
  // pam3_sub_sys_TEA_f1
  output logic           pam3_sub_sys_TEA_f1_activity,                          // Upcoming activity indicator
  output logic           pam3_sub_sys_TEA_f1_req,                               // Flit transfer request
  output logic           pam3_sub_sys_TEA_f1_sop,                               // Start of packet indicator
  output logic           pam3_sub_sys_TEA_f1_eop,                               // End of packet indicator
  output logic    [59:0] pam3_sub_sys_TEA_f1_flitdata,                          // Flit data
  input  wire            pam3_sub_sys_TEA_f1_ready,                             // Flit transfer ready
  // pam3_sub_sys_TEA_r0
  input  wire            pam3_sub_sys_TEA_r0_activity,                          // Upcoming activity indicator
  input  wire            pam3_sub_sys_TEA_r0_req,                               // Flit transfer request
  input  wire            pam3_sub_sys_TEA_r0_sop,                               // Start of packet indicator
  input  wire            pam3_sub_sys_TEA_r0_eop,                               // End of packet indicator
  input  wire     [33:0] pam3_sub_sys_TEA_r0_flitdata,                          // Flit data
  output logic           pam3_sub_sys_TEA_r0_ready,                             // Flit transfer ready
  // pam3_sub_sys_TEA_r1
  input  wire            pam3_sub_sys_TEA_r1_activity,                          // Upcoming activity indicator
  input  wire            pam3_sub_sys_TEA_r1_req,                               // Flit transfer request
  input  wire            pam3_sub_sys_TEA_r1_sop,                               // Start of packet indicator
  input  wire            pam3_sub_sys_TEA_r1_eop,                               // End of packet indicator
  input  wire     [23:0] pam3_sub_sys_TEA_r1_flitdata,                          // Flit data
  output logic           pam3_sub_sys_TEA_r1_ready,                             // Flit transfer ready
  // usb4_phy_TEA_f0
  output logic           usb4_phy_TEA_f0_activity,                              // Upcoming activity indicator
  output logic           usb4_phy_TEA_f0_req,                                   // Flit transfer request
  output logic           usb4_phy_TEA_f0_sop,                                   // Start of packet indicator
  output logic           usb4_phy_TEA_f0_eop,                                   // End of packet indicator
  output logic    [35:0] usb4_phy_TEA_f0_flitdata,                              // Flit data
  input  wire            usb4_phy_TEA_f0_ready,                                 // Flit transfer ready
  // usb4_phy_TEA_f1
  output logic           usb4_phy_TEA_f1_activity,                              // Upcoming activity indicator
  output logic           usb4_phy_TEA_f1_req,                                   // Flit transfer request
  output logic           usb4_phy_TEA_f1_sop,                                   // Start of packet indicator
  output logic           usb4_phy_TEA_f1_eop,                                   // End of packet indicator
  output logic    [59:0] usb4_phy_TEA_f1_flitdata,                              // Flit data
  input  wire            usb4_phy_TEA_f1_ready,                                 // Flit transfer ready
  // usb4_phy_TEA_r0
  input  wire            usb4_phy_TEA_r0_activity,                              // Upcoming activity indicator
  input  wire            usb4_phy_TEA_r0_req,                                   // Flit transfer request
  input  wire            usb4_phy_TEA_r0_sop,                                   // Start of packet indicator
  input  wire            usb4_phy_TEA_r0_eop,                                   // End of packet indicator
  input  wire     [33:0] usb4_phy_TEA_r0_flitdata,                              // Flit data
  output logic           usb4_phy_TEA_r0_ready,                                 // Flit transfer ready
  // usb4_phy_TEA_r1
  input  wire            usb4_phy_TEA_r1_activity,                              // Upcoming activity indicator
  input  wire            usb4_phy_TEA_r1_req,                                   // Flit transfer request
  input  wire            usb4_phy_TEA_r1_sop,                                   // Start of packet indicator
  input  wire            usb4_phy_TEA_r1_eop,                                   // End of packet indicator
  input  wire     [23:0] usb4_phy_TEA_r1_flitdata,                              // Flit data
  output logic           usb4_phy_TEA_r1_ready,                                 // Flit transfer ready
  // pam3_xcvr_TEA_f0
  output logic           pam3_xcvr_TEA_f0_activity,                             // Upcoming activity indicator
  output logic           pam3_xcvr_TEA_f0_req,                                  // Flit transfer request
  output logic           pam3_xcvr_TEA_f0_sop,                                  // Start of packet indicator
  output logic           pam3_xcvr_TEA_f0_eop,                                  // End of packet indicator
  output logic    [35:0] pam3_xcvr_TEA_f0_flitdata,                             // Flit data
  input  wire            pam3_xcvr_TEA_f0_ready,                                // Flit transfer ready
  // pam3_xcvr_TEA_f1
  output logic           pam3_xcvr_TEA_f1_activity,                             // Upcoming activity indicator
  output logic           pam3_xcvr_TEA_f1_req,                                  // Flit transfer request
  output logic           pam3_xcvr_TEA_f1_sop,                                  // Start of packet indicator
  output logic           pam3_xcvr_TEA_f1_eop,                                  // End of packet indicator
  output logic    [59:0] pam3_xcvr_TEA_f1_flitdata,                             // Flit data
  input  wire            pam3_xcvr_TEA_f1_ready,                                // Flit transfer ready
  // pam3_xcvr_TEA_r0
  input  wire            pam3_xcvr_TEA_r0_activity,                             // Upcoming activity indicator
  input  wire            pam3_xcvr_TEA_r0_req,                                  // Flit transfer request
  input  wire            pam3_xcvr_TEA_r0_sop,                                  // Start of packet indicator
  input  wire            pam3_xcvr_TEA_r0_eop,                                  // End of packet indicator
  input  wire     [33:0] pam3_xcvr_TEA_r0_flitdata,                             // Flit data
  output logic           pam3_xcvr_TEA_r0_ready,                                // Flit transfer ready
  // pam3_xcvr_TEA_r1
  input  wire            pam3_xcvr_TEA_r1_activity,                             // Upcoming activity indicator
  input  wire            pam3_xcvr_TEA_r1_req,                                  // Flit transfer request
  input  wire            pam3_xcvr_TEA_r1_sop,                                  // Start of packet indicator
  input  wire            pam3_xcvr_TEA_r1_eop,                                  // End of packet indicator
  input  wire     [23:0] pam3_xcvr_TEA_r1_flitdata,                             // Flit data
  output logic           pam3_xcvr_TEA_r1_ready                                 // Flit transfer ready
);

logic           trigger;
logic           f0_i0_sop;
logic           f0_i0_eop;
logic     [3:0] f0_i0_qos_nxt;
logic     [3:0] f0_i0_qos;
logic    [35:0] f0_i0_flitdata;
logic           f0_i0_t4_activity;
logic           f0_i0_t4_req_nxt;
logic           f0_i0_t4_req;
logic           f0_i0_t4_ready;
logic           f0_i0_t2_activity;
logic           f0_i0_t2_req_nxt;
logic           f0_i0_t2_req;
logic           f0_i0_t2_ready;
logic           f0_i0_t1_activity;
logic           f0_i0_t1_req_nxt;
logic           f0_i0_t1_req;
logic           f0_i0_t1_ready;
logic           f0_i0_t0_activity;
logic           f0_i0_t0_req_nxt;
logic           f0_i0_t0_req;
logic           f0_i0_t0_ready;
logic           f0_i0_t5_activity;
logic           f0_i0_t5_req_nxt;
logic           f0_i0_t5_req;
logic           f0_i0_t5_ready;
logic           f0_i0_t3_activity;
logic           f0_i0_t3_req_nxt;
logic           f0_i0_t3_req;
logic           f0_i0_t3_ready;
logic           f0_i0_t1000_activity;
logic           f0_i0_t1000_req_nxt;
logic           f0_i0_t1000_req;
logic           f0_i0_t1000_ready;
logic           f1_i0_sop;
logic           f1_i0_eop;
logic     [3:0] f1_i0_qos_nxt;
logic     [3:0] f1_i0_qos;
logic    [59:0] f1_i0_flitdata;
logic           f1_i0_t4_activity;
logic           f1_i0_t4_req_nxt;
logic           f1_i0_t4_req;
logic           f1_i0_t4_ready;
logic           f1_i0_t2_activity;
logic           f1_i0_t2_req_nxt;
logic           f1_i0_t2_req;
logic           f1_i0_t2_ready;
logic           f1_i0_t1_activity;
logic           f1_i0_t1_req_nxt;
logic           f1_i0_t1_req;
logic           f1_i0_t1_ready;
logic           f1_i0_t0_activity;
logic           f1_i0_t0_req_nxt;
logic           f1_i0_t0_req;
logic           f1_i0_t0_ready;
logic           f1_i0_t5_activity;
logic           f1_i0_t5_req_nxt;
logic           f1_i0_t5_req;
logic           f1_i0_t5_ready;
logic           f1_i0_t3_activity;
logic           f1_i0_t3_req_nxt;
logic           f1_i0_t3_req;
logic           f1_i0_t3_ready;
logic           f1_i0_t1000_activity;
logic           f1_i0_t1000_req_nxt;
logic           f1_i0_t1000_req;
logic           f1_i0_t1000_ready;
logic           f0_i1_sop;
logic           f0_i1_eop;
logic     [3:0] f0_i1_qos_nxt;
logic     [3:0] f0_i1_qos;
logic    [35:0] f0_i1_flitdata;
logic           f0_i1_t4_activity;
logic           f0_i1_t4_req_nxt;
logic           f0_i1_t4_req;
logic           f0_i1_t4_ready;
logic           f0_i1_t2_activity;
logic           f0_i1_t2_req_nxt;
logic           f0_i1_t2_req;
logic           f0_i1_t2_ready;
logic           f0_i1_t1_activity;
logic           f0_i1_t1_req_nxt;
logic           f0_i1_t1_req;
logic           f0_i1_t1_ready;
logic           f0_i1_t0_activity;
logic           f0_i1_t0_req_nxt;
logic           f0_i1_t0_req;
logic           f0_i1_t0_ready;
logic           f0_i1_t5_activity;
logic           f0_i1_t5_req_nxt;
logic           f0_i1_t5_req;
logic           f0_i1_t5_ready;
logic           f0_i1_t3_activity;
logic           f0_i1_t3_req_nxt;
logic           f0_i1_t3_req;
logic           f0_i1_t3_ready;
logic           f0_i1_t1000_activity;
logic           f0_i1_t1000_req_nxt;
logic           f0_i1_t1000_req;
logic           f0_i1_t1000_ready;
logic           f1_i1_sop;
logic           f1_i1_eop;
logic     [3:0] f1_i1_qos_nxt;
logic     [3:0] f1_i1_qos;
logic    [59:0] f1_i1_flitdata;
logic           f1_i1_t4_activity;
logic           f1_i1_t4_req_nxt;
logic           f1_i1_t4_req;
logic           f1_i1_t4_ready;
logic           f1_i1_t2_activity;
logic           f1_i1_t2_req_nxt;
logic           f1_i1_t2_req;
logic           f1_i1_t2_ready;
logic           f1_i1_t1_activity;
logic           f1_i1_t1_req_nxt;
logic           f1_i1_t1_req;
logic           f1_i1_t1_ready;
logic           f1_i1_t0_activity;
logic           f1_i1_t0_req_nxt;
logic           f1_i1_t0_req;
logic           f1_i1_t0_ready;
logic           f1_i1_t5_activity;
logic           f1_i1_t5_req_nxt;
logic           f1_i1_t5_req;
logic           f1_i1_t5_ready;
logic           f1_i1_t3_activity;
logic           f1_i1_t3_req_nxt;
logic           f1_i1_t3_req;
logic           f1_i1_t3_ready;
logic           f1_i1_t1000_activity;
logic           f1_i1_t1000_req_nxt;
logic           f1_i1_t1000_req;
logic           f1_i1_t1000_ready;
logic           r0_t0_sop;
logic           r0_t0_eop;
logic     [3:0] r0_t0_qos_nxt;
logic     [3:0] r0_t0_qos;
logic    [33:0] r0_t0_flitdata;
logic           r0_t0_i0_activity;
logic           r0_t0_i0_req_nxt;
logic           r0_t0_i0_req;
logic           r0_t0_i0_ready;
logic           r0_t0_i1_activity;
logic           r0_t0_i1_req_nxt;
logic           r0_t0_i1_req;
logic           r0_t0_i1_ready;
logic           r1_t0_sop;
logic           r1_t0_eop;
logic     [3:0] r1_t0_qos_nxt;
logic     [3:0] r1_t0_qos;
logic    [23:0] r1_t0_flitdata;
logic           r1_t0_i0_activity;
logic           r1_t0_i0_req_nxt;
logic           r1_t0_i0_req;
logic           r1_t0_i0_ready;
logic           r1_t0_i1_activity;
logic           r1_t0_i1_req_nxt;
logic           r1_t0_i1_req;
logic           r1_t0_i1_ready;
logic           r0_t1_sop;
logic           r0_t1_eop;
logic     [3:0] r0_t1_qos_nxt;
logic     [3:0] r0_t1_qos;
logic    [33:0] r0_t1_flitdata;
logic           r0_t1_i0_activity;
logic           r0_t1_i0_req_nxt;
logic           r0_t1_i0_req;
logic           r0_t1_i0_ready;
logic           r0_t1_i1_activity;
logic           r0_t1_i1_req_nxt;
logic           r0_t1_i1_req;
logic           r0_t1_i1_ready;
logic           r1_t1_sop;
logic           r1_t1_eop;
logic     [3:0] r1_t1_qos_nxt;
logic     [3:0] r1_t1_qos;
logic    [23:0] r1_t1_flitdata;
logic           r1_t1_i0_activity;
logic           r1_t1_i0_req_nxt;
logic           r1_t1_i0_req;
logic           r1_t1_i0_ready;
logic           r1_t1_i1_activity;
logic           r1_t1_i1_req_nxt;
logic           r1_t1_i1_req;
logic           r1_t1_i1_ready;
logic           r0_t2_sop;
logic           r0_t2_eop;
logic     [3:0] r0_t2_qos_nxt;
logic     [3:0] r0_t2_qos;
logic    [33:0] r0_t2_flitdata;
logic           r0_t2_i0_activity;
logic           r0_t2_i0_req_nxt;
logic           r0_t2_i0_req;
logic           r0_t2_i0_ready;
logic           r0_t2_i1_activity;
logic           r0_t2_i1_req_nxt;
logic           r0_t2_i1_req;
logic           r0_t2_i1_ready;
logic           r1_t2_sop;
logic           r1_t2_eop;
logic     [3:0] r1_t2_qos_nxt;
logic     [3:0] r1_t2_qos;
logic    [23:0] r1_t2_flitdata;
logic           r1_t2_i0_activity;
logic           r1_t2_i0_req_nxt;
logic           r1_t2_i0_req;
logic           r1_t2_i0_ready;
logic           r1_t2_i1_activity;
logic           r1_t2_i1_req_nxt;
logic           r1_t2_i1_req;
logic           r1_t2_i1_ready;
logic           r0_t3_sop;
logic           r0_t3_eop;
logic     [3:0] r0_t3_qos_nxt;
logic     [3:0] r0_t3_qos;
logic    [33:0] r0_t3_flitdata;
logic           r0_t3_i0_activity;
logic           r0_t3_i0_req_nxt;
logic           r0_t3_i0_req;
logic           r0_t3_i0_ready;
logic           r0_t3_i1_activity;
logic           r0_t3_i1_req_nxt;
logic           r0_t3_i1_req;
logic           r0_t3_i1_ready;
logic           r1_t3_sop;
logic           r1_t3_eop;
logic     [3:0] r1_t3_qos_nxt;
logic     [3:0] r1_t3_qos;
logic    [23:0] r1_t3_flitdata;
logic           r1_t3_i0_activity;
logic           r1_t3_i0_req_nxt;
logic           r1_t3_i0_req;
logic           r1_t3_i0_ready;
logic           r1_t3_i1_activity;
logic           r1_t3_i1_req_nxt;
logic           r1_t3_i1_req;
logic           r1_t3_i1_ready;
logic           r0_t4_sop;
logic           r0_t4_eop;
logic     [3:0] r0_t4_qos_nxt;
logic     [3:0] r0_t4_qos;
logic    [33:0] r0_t4_flitdata;
logic           r0_t4_i0_activity;
logic           r0_t4_i0_req_nxt;
logic           r0_t4_i0_req;
logic           r0_t4_i0_ready;
logic           r0_t4_i1_activity;
logic           r0_t4_i1_req_nxt;
logic           r0_t4_i1_req;
logic           r0_t4_i1_ready;
logic           r1_t4_sop;
logic           r1_t4_eop;
logic     [3:0] r1_t4_qos_nxt;
logic     [3:0] r1_t4_qos;
logic    [23:0] r1_t4_flitdata;
logic           r1_t4_i0_activity;
logic           r1_t4_i0_req_nxt;
logic           r1_t4_i0_req;
logic           r1_t4_i0_ready;
logic           r1_t4_i1_activity;
logic           r1_t4_i1_req_nxt;
logic           r1_t4_i1_req;
logic           r1_t4_i1_ready;
logic           r0_t5_sop;
logic           r0_t5_eop;
logic     [3:0] r0_t5_qos_nxt;
logic     [3:0] r0_t5_qos;
logic    [33:0] r0_t5_flitdata;
logic           r0_t5_i0_activity;
logic           r0_t5_i0_req_nxt;
logic           r0_t5_i0_req;
logic           r0_t5_i0_ready;
logic           r0_t5_i1_activity;
logic           r0_t5_i1_req_nxt;
logic           r0_t5_i1_req;
logic           r0_t5_i1_ready;
logic           r1_t5_sop;
logic           r1_t5_eop;
logic     [3:0] r1_t5_qos_nxt;
logic     [3:0] r1_t5_qos;
logic    [23:0] r1_t5_flitdata;
logic           r1_t5_i0_activity;
logic           r1_t5_i0_req_nxt;
logic           r1_t5_i0_req;
logic           r1_t5_i0_ready;
logic           r1_t5_i1_activity;
logic           r1_t5_i1_req_nxt;
logic           r1_t5_i1_req;
logic           r1_t5_i1_ready;
logic           r0_t1000_sop;
logic           r0_t1000_eop;
logic     [3:0] r0_t1000_qos_nxt;
logic     [3:0] r0_t1000_qos;
logic    [33:0] r0_t1000_flitdata;
logic           r0_t1000_i0_activity;
logic           r0_t1000_i0_req_nxt;
logic           r0_t1000_i0_req;
logic           r0_t1000_i0_ready;
logic           r0_t1000_i1_activity;
logic           r0_t1000_i1_req_nxt;
logic           r0_t1000_i1_req;
logic           r0_t1000_i1_ready;
logic           r1_t1000_sop;
logic           r1_t1000_eop;
logic     [3:0] r1_t1000_qos_nxt;
logic     [3:0] r1_t1000_qos;
logic    [23:0] r1_t1000_flitdata;
logic           r1_t1000_i0_activity;
logic           r1_t1000_i0_req_nxt;
logic           r1_t1000_i0_req;
logic           r1_t1000_i0_ready;
logic           r1_t1000_i1_activity;
logic           r1_t1000_i1_req_nxt;
logic           r1_t1000_i1_req;
logic           r1_t1000_i1_ready;
logic           regWReq;
logic     [9:0] regWAddr;
logic    [31:0] regWData;
logic     [3:0] regWEn;
logic           regRReq;
logic     [9:0] regRAddr;
logic    [31:0] regRData;
logic           t1000_f0_activity;                                              // Upcoming activity indicator
logic           t1000_f0_req;                                                   // Flit transfer request
logic           t1000_f0_sop;                                                   // Start of packet indicator
logic           t1000_f0_eop;                                                   // End of packet indicator
logic    [35:0] t1000_f0_flitdata;                                              // Flit data
logic           t1000_f0_ready;                                                 // Flit transfer ready
logic           t1000_f1_activity;                                              // Upcoming activity indicator
logic           t1000_f1_req;                                                   // Flit transfer request
logic           t1000_f1_sop;                                                   // Start of packet indicator
logic           t1000_f1_eop;                                                   // End of packet indicator
logic    [59:0] t1000_f1_flitdata;                                              // Flit data
logic           t1000_f1_ready;                                                 // Flit transfer ready
logic           t1000_r0_activity;                                              // Upcoming activity indicator
logic           t1000_r0_req;                                                   // Flit transfer request
logic           t1000_r0_sop;                                                   // Start of packet indicator
logic           t1000_r0_eop;                                                   // End of packet indicator
logic    [33:0] t1000_r0_flitdata;                                              // Flit data
logic           t1000_r0_ready;                                                 // Flit transfer ready
logic           t1000_r1_activity;                                              // Upcoming activity indicator
logic           t1000_r1_req;                                                   // Flit transfer request
logic           t1000_r1_sop;                                                   // Start of packet indicator
logic           t1000_r1_eop;                                                   // End of packet indicator
logic    [23:0] t1000_r1_flitdata;                                              // Flit data
logic           t1000_r1_ready;                                                 // Flit transfer ready
logic           frst_n;                                                         // Output reset for async flops
logic           lrst_n;                                                         // Output reset for everything else
logic     [0:0] t1000_f0_srcIdx;
logic     [0:0] t1000_f1_srcIdx;
logic     [0:0] t1000_r0_dstIdx;
logic     [0:0] t1000_r1_dstIdx;
logic    [47:0] monCnt;
logic    [47:0] monCnt_nxt;
logic     [0:0] monCnt_en;
logic           monRunning;
logic     [0:0] monSet;
logic     [0:0] monSet_nxt;
logic     [0:0] monSet_en;
logic     [0:0] monUpd;
logic     [0:0] monUpd_nxt;
logic     [0:0] monUpd_en;
logic     [1:0] monMode;
logic     [1:0] monMode_nxt;
logic     [0:0] monMode_en;
logic     [3:0] regMSB;
logic           newMode;
logic    [31:0] regData [3:0];
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
usb4_tc_noc_rtr0_rstS rstS (
  .clk(clk),                                                                    // i:1
  .rawReset(rst_n),                                                             // i:1
  .flopReset(frst_n),                                                           // o:1
  .logicReset(lrst_n)                                                           // o:1
);
// ============================================================================
// Synchronize any isolation link pins
// ============================================================================
// ============================================================================
// ============================================================================
// Initiator Interfaces
// ============================================================================
// ============================================================================
// ============================================================================
// Initiator Port 0 Forward Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Initiator Port 0 Forward Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_f0_dec apb_mstr_f0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .trigger(trigger),                                                            // i:1
  .ini_activity(apb_mstr_f0_activity),                                          // i:1
  .ini_req(apb_mstr_f0_req),                                                    // i:1
  .ini_sop(apb_mstr_f0_sop),                                                    // i:1
  .ini_eop(apb_mstr_f0_eop),                                                    // i:1
  .ini_flitdata(apb_mstr_f0_flitdata),                                          // i:36
  .ini_ready(apb_mstr_f0_ready),                                                // o:1
  .f0_i0_sop(f0_i0_sop),                                                        // o:1
  .f0_i0_eop(f0_i0_eop),                                                        // o:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // o:4
  .f0_i0_qos(f0_i0_qos),                                                        // o:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // o:36
  .f0_i0_t4_activity(f0_i0_t4_activity),                                        // o:1
  .f0_i0_t4_req_nxt(f0_i0_t4_req_nxt),                                          // o:1
  .f0_i0_t4_req(f0_i0_t4_req),                                                  // o:1
  .f0_i0_t4_ready(f0_i0_t4_ready),                                              // i:1
  .f0_i0_t2_activity(f0_i0_t2_activity),                                        // o:1
  .f0_i0_t2_req_nxt(f0_i0_t2_req_nxt),                                          // o:1
  .f0_i0_t2_req(f0_i0_t2_req),                                                  // o:1
  .f0_i0_t2_ready(f0_i0_t2_ready),                                              // i:1
  .f0_i0_t1_activity(f0_i0_t1_activity),                                        // o:1
  .f0_i0_t1_req_nxt(f0_i0_t1_req_nxt),                                          // o:1
  .f0_i0_t1_req(f0_i0_t1_req),                                                  // o:1
  .f0_i0_t1_ready(f0_i0_t1_ready),                                              // i:1
  .f0_i0_t0_activity(f0_i0_t0_activity),                                        // o:1
  .f0_i0_t0_req_nxt(f0_i0_t0_req_nxt),                                          // o:1
  .f0_i0_t0_req(f0_i0_t0_req),                                                  // o:1
  .f0_i0_t0_ready(f0_i0_t0_ready),                                              // i:1
  .f0_i0_t5_activity(f0_i0_t5_activity),                                        // o:1
  .f0_i0_t5_req_nxt(f0_i0_t5_req_nxt),                                          // o:1
  .f0_i0_t5_req(f0_i0_t5_req),                                                  // o:1
  .f0_i0_t5_ready(f0_i0_t5_ready),                                              // i:1
  .f0_i0_t3_activity(f0_i0_t3_activity),                                        // o:1
  .f0_i0_t3_req_nxt(f0_i0_t3_req_nxt),                                          // o:1
  .f0_i0_t3_req(f0_i0_t3_req),                                                  // o:1
  .f0_i0_t3_ready(f0_i0_t3_ready),                                              // i:1
  .f0_i0_t1000_activity(f0_i0_t1000_activity),                                  // o:1
  .f0_i0_t1000_req_nxt(f0_i0_t1000_req_nxt),                                    // o:1
  .f0_i0_t1000_req(f0_i0_t1000_req),                                            // o:1
  .f0_i0_t1000_ready(f0_i0_t1000_ready)                                         // i:1
);
// ============================================================================
// Initiator Port 0 Forward Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Initiator Port 0 Forward Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_f1_dec apb_mstr_f1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .trigger(trigger),                                                            // i:1
  .ini_activity(apb_mstr_f1_activity),                                          // i:1
  .ini_req(apb_mstr_f1_req),                                                    // i:1
  .ini_sop(apb_mstr_f1_sop),                                                    // i:1
  .ini_eop(apb_mstr_f1_eop),                                                    // i:1
  .ini_flitdata(apb_mstr_f1_flitdata),                                          // i:60
  .ini_ready(apb_mstr_f1_ready),                                                // o:1
  .f1_i0_sop(f1_i0_sop),                                                        // o:1
  .f1_i0_eop(f1_i0_eop),                                                        // o:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // o:4
  .f1_i0_qos(f1_i0_qos),                                                        // o:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // o:60
  .f1_i0_t4_activity(f1_i0_t4_activity),                                        // o:1
  .f1_i0_t4_req_nxt(f1_i0_t4_req_nxt),                                          // o:1
  .f1_i0_t4_req(f1_i0_t4_req),                                                  // o:1
  .f1_i0_t4_ready(f1_i0_t4_ready),                                              // i:1
  .f1_i0_t2_activity(f1_i0_t2_activity),                                        // o:1
  .f1_i0_t2_req_nxt(f1_i0_t2_req_nxt),                                          // o:1
  .f1_i0_t2_req(f1_i0_t2_req),                                                  // o:1
  .f1_i0_t2_ready(f1_i0_t2_ready),                                              // i:1
  .f1_i0_t1_activity(f1_i0_t1_activity),                                        // o:1
  .f1_i0_t1_req_nxt(f1_i0_t1_req_nxt),                                          // o:1
  .f1_i0_t1_req(f1_i0_t1_req),                                                  // o:1
  .f1_i0_t1_ready(f1_i0_t1_ready),                                              // i:1
  .f1_i0_t0_activity(f1_i0_t0_activity),                                        // o:1
  .f1_i0_t0_req_nxt(f1_i0_t0_req_nxt),                                          // o:1
  .f1_i0_t0_req(f1_i0_t0_req),                                                  // o:1
  .f1_i0_t0_ready(f1_i0_t0_ready),                                              // i:1
  .f1_i0_t5_activity(f1_i0_t5_activity),                                        // o:1
  .f1_i0_t5_req_nxt(f1_i0_t5_req_nxt),                                          // o:1
  .f1_i0_t5_req(f1_i0_t5_req),                                                  // o:1
  .f1_i0_t5_ready(f1_i0_t5_ready),                                              // i:1
  .f1_i0_t3_activity(f1_i0_t3_activity),                                        // o:1
  .f1_i0_t3_req_nxt(f1_i0_t3_req_nxt),                                          // o:1
  .f1_i0_t3_req(f1_i0_t3_req),                                                  // o:1
  .f1_i0_t3_ready(f1_i0_t3_ready),                                              // i:1
  .f1_i0_t1000_activity(f1_i0_t1000_activity),                                  // o:1
  .f1_i0_t1000_req_nxt(f1_i0_t1000_req_nxt),                                    // o:1
  .f1_i0_t1000_req(f1_i0_t1000_req),                                            // o:1
  .f1_i0_t1000_ready(f1_i0_t1000_ready)                                         // i:1
);
// ============================================================================
// Initiator Port 0 Reverse Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Initiator Port 0 Reverse Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_r0_arb apb_mstr_r0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .r0_t4_sop(r0_t4_sop),                                                        // i:1
  .r0_t4_eop(r0_t4_eop),                                                        // i:1
  .r0_t4_qos_nxt(r0_t4_qos_nxt),                                                // i:4
  .r0_t4_qos(r0_t4_qos),                                                        // i:4
  .r0_t4_flitdata(r0_t4_flitdata),                                              // i:34
  .r0_t4_i0_activity(r0_t4_i0_activity),                                        // i:1
  .r0_t4_i0_req_nxt(r0_t4_i0_req_nxt),                                          // i:1
  .r0_t4_i0_req(r0_t4_i0_req),                                                  // i:1
  .r0_t4_i0_ready(r0_t4_i0_ready),                                              // o:1
  .r0_t2_sop(r0_t2_sop),                                                        // i:1
  .r0_t2_eop(r0_t2_eop),                                                        // i:1
  .r0_t2_qos_nxt(r0_t2_qos_nxt),                                                // i:4
  .r0_t2_qos(r0_t2_qos),                                                        // i:4
  .r0_t2_flitdata(r0_t2_flitdata),                                              // i:34
  .r0_t2_i0_activity(r0_t2_i0_activity),                                        // i:1
  .r0_t2_i0_req_nxt(r0_t2_i0_req_nxt),                                          // i:1
  .r0_t2_i0_req(r0_t2_i0_req),                                                  // i:1
  .r0_t2_i0_ready(r0_t2_i0_ready),                                              // o:1
  .r0_t1_sop(r0_t1_sop),                                                        // i:1
  .r0_t1_eop(r0_t1_eop),                                                        // i:1
  .r0_t1_qos_nxt(r0_t1_qos_nxt),                                                // i:4
  .r0_t1_qos(r0_t1_qos),                                                        // i:4
  .r0_t1_flitdata(r0_t1_flitdata),                                              // i:34
  .r0_t1_i0_activity(r0_t1_i0_activity),                                        // i:1
  .r0_t1_i0_req_nxt(r0_t1_i0_req_nxt),                                          // i:1
  .r0_t1_i0_req(r0_t1_i0_req),                                                  // i:1
  .r0_t1_i0_ready(r0_t1_i0_ready),                                              // o:1
  .r0_t0_sop(r0_t0_sop),                                                        // i:1
  .r0_t0_eop(r0_t0_eop),                                                        // i:1
  .r0_t0_qos_nxt(r0_t0_qos_nxt),                                                // i:4
  .r0_t0_qos(r0_t0_qos),                                                        // i:4
  .r0_t0_flitdata(r0_t0_flitdata),                                              // i:34
  .r0_t0_i0_activity(r0_t0_i0_activity),                                        // i:1
  .r0_t0_i0_req_nxt(r0_t0_i0_req_nxt),                                          // i:1
  .r0_t0_i0_req(r0_t0_i0_req),                                                  // i:1
  .r0_t0_i0_ready(r0_t0_i0_ready),                                              // o:1
  .r0_t5_sop(r0_t5_sop),                                                        // i:1
  .r0_t5_eop(r0_t5_eop),                                                        // i:1
  .r0_t5_qos_nxt(r0_t5_qos_nxt),                                                // i:4
  .r0_t5_qos(r0_t5_qos),                                                        // i:4
  .r0_t5_flitdata(r0_t5_flitdata),                                              // i:34
  .r0_t5_i0_activity(r0_t5_i0_activity),                                        // i:1
  .r0_t5_i0_req_nxt(r0_t5_i0_req_nxt),                                          // i:1
  .r0_t5_i0_req(r0_t5_i0_req),                                                  // i:1
  .r0_t5_i0_ready(r0_t5_i0_ready),                                              // o:1
  .r0_t3_sop(r0_t3_sop),                                                        // i:1
  .r0_t3_eop(r0_t3_eop),                                                        // i:1
  .r0_t3_qos_nxt(r0_t3_qos_nxt),                                                // i:4
  .r0_t3_qos(r0_t3_qos),                                                        // i:4
  .r0_t3_flitdata(r0_t3_flitdata),                                              // i:34
  .r0_t3_i0_activity(r0_t3_i0_activity),                                        // i:1
  .r0_t3_i0_req_nxt(r0_t3_i0_req_nxt),                                          // i:1
  .r0_t3_i0_req(r0_t3_i0_req),                                                  // i:1
  .r0_t3_i0_ready(r0_t3_i0_ready),                                              // o:1
  .r0_t1000_sop(r0_t1000_sop),                                                  // i:1
  .r0_t1000_eop(r0_t1000_eop),                                                  // i:1
  .r0_t1000_qos_nxt(r0_t1000_qos_nxt),                                          // i:4
  .r0_t1000_qos(r0_t1000_qos),                                                  // i:4
  .r0_t1000_flitdata(r0_t1000_flitdata),                                        // i:34
  .r0_t1000_i0_activity(r0_t1000_i0_activity),                                  // i:1
  .r0_t1000_i0_req_nxt(r0_t1000_i0_req_nxt),                                    // i:1
  .r0_t1000_i0_req(r0_t1000_i0_req),                                            // i:1
  .r0_t1000_i0_ready(r0_t1000_i0_ready),                                        // o:1
  .tgt_activity(apb_mstr_r0_activity),                                          // o:1
  .tgt_req(apb_mstr_r0_req),                                                    // o:1
  .tgt_sop(apb_mstr_r0_sop),                                                    // o:1
  .tgt_eop(apb_mstr_r0_eop),                                                    // o:1
  .tgt_flitdata(apb_mstr_r0_flitdata),                                          // o:34
  .tgt_ready(apb_mstr_r0_ready)                                                 // i:1
);
// ============================================================================
// Initiator Port 0 Reverse Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Initiator Port 0 Reverse Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_r1_arb apb_mstr_r1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .r1_t4_sop(r1_t4_sop),                                                        // i:1
  .r1_t4_eop(r1_t4_eop),                                                        // i:1
  .r1_t4_qos_nxt(r1_t4_qos_nxt),                                                // i:4
  .r1_t4_qos(r1_t4_qos),                                                        // i:4
  .r1_t4_flitdata(r1_t4_flitdata),                                              // i:24
  .r1_t4_i0_activity(r1_t4_i0_activity),                                        // i:1
  .r1_t4_i0_req_nxt(r1_t4_i0_req_nxt),                                          // i:1
  .r1_t4_i0_req(r1_t4_i0_req),                                                  // i:1
  .r1_t4_i0_ready(r1_t4_i0_ready),                                              // o:1
  .r1_t2_sop(r1_t2_sop),                                                        // i:1
  .r1_t2_eop(r1_t2_eop),                                                        // i:1
  .r1_t2_qos_nxt(r1_t2_qos_nxt),                                                // i:4
  .r1_t2_qos(r1_t2_qos),                                                        // i:4
  .r1_t2_flitdata(r1_t2_flitdata),                                              // i:24
  .r1_t2_i0_activity(r1_t2_i0_activity),                                        // i:1
  .r1_t2_i0_req_nxt(r1_t2_i0_req_nxt),                                          // i:1
  .r1_t2_i0_req(r1_t2_i0_req),                                                  // i:1
  .r1_t2_i0_ready(r1_t2_i0_ready),                                              // o:1
  .r1_t1_sop(r1_t1_sop),                                                        // i:1
  .r1_t1_eop(r1_t1_eop),                                                        // i:1
  .r1_t1_qos_nxt(r1_t1_qos_nxt),                                                // i:4
  .r1_t1_qos(r1_t1_qos),                                                        // i:4
  .r1_t1_flitdata(r1_t1_flitdata),                                              // i:24
  .r1_t1_i0_activity(r1_t1_i0_activity),                                        // i:1
  .r1_t1_i0_req_nxt(r1_t1_i0_req_nxt),                                          // i:1
  .r1_t1_i0_req(r1_t1_i0_req),                                                  // i:1
  .r1_t1_i0_ready(r1_t1_i0_ready),                                              // o:1
  .r1_t0_sop(r1_t0_sop),                                                        // i:1
  .r1_t0_eop(r1_t0_eop),                                                        // i:1
  .r1_t0_qos_nxt(r1_t0_qos_nxt),                                                // i:4
  .r1_t0_qos(r1_t0_qos),                                                        // i:4
  .r1_t0_flitdata(r1_t0_flitdata),                                              // i:24
  .r1_t0_i0_activity(r1_t0_i0_activity),                                        // i:1
  .r1_t0_i0_req_nxt(r1_t0_i0_req_nxt),                                          // i:1
  .r1_t0_i0_req(r1_t0_i0_req),                                                  // i:1
  .r1_t0_i0_ready(r1_t0_i0_ready),                                              // o:1
  .r1_t5_sop(r1_t5_sop),                                                        // i:1
  .r1_t5_eop(r1_t5_eop),                                                        // i:1
  .r1_t5_qos_nxt(r1_t5_qos_nxt),                                                // i:4
  .r1_t5_qos(r1_t5_qos),                                                        // i:4
  .r1_t5_flitdata(r1_t5_flitdata),                                              // i:24
  .r1_t5_i0_activity(r1_t5_i0_activity),                                        // i:1
  .r1_t5_i0_req_nxt(r1_t5_i0_req_nxt),                                          // i:1
  .r1_t5_i0_req(r1_t5_i0_req),                                                  // i:1
  .r1_t5_i0_ready(r1_t5_i0_ready),                                              // o:1
  .r1_t3_sop(r1_t3_sop),                                                        // i:1
  .r1_t3_eop(r1_t3_eop),                                                        // i:1
  .r1_t3_qos_nxt(r1_t3_qos_nxt),                                                // i:4
  .r1_t3_qos(r1_t3_qos),                                                        // i:4
  .r1_t3_flitdata(r1_t3_flitdata),                                              // i:24
  .r1_t3_i0_activity(r1_t3_i0_activity),                                        // i:1
  .r1_t3_i0_req_nxt(r1_t3_i0_req_nxt),                                          // i:1
  .r1_t3_i0_req(r1_t3_i0_req),                                                  // i:1
  .r1_t3_i0_ready(r1_t3_i0_ready),                                              // o:1
  .r1_t1000_sop(r1_t1000_sop),                                                  // i:1
  .r1_t1000_eop(r1_t1000_eop),                                                  // i:1
  .r1_t1000_qos_nxt(r1_t1000_qos_nxt),                                          // i:4
  .r1_t1000_qos(r1_t1000_qos),                                                  // i:4
  .r1_t1000_flitdata(r1_t1000_flitdata),                                        // i:24
  .r1_t1000_i0_activity(r1_t1000_i0_activity),                                  // i:1
  .r1_t1000_i0_req_nxt(r1_t1000_i0_req_nxt),                                    // i:1
  .r1_t1000_i0_req(r1_t1000_i0_req),                                            // i:1
  .r1_t1000_i0_ready(r1_t1000_i0_ready),                                        // o:1
  .tgt_activity(apb_mstr_r1_activity),                                          // o:1
  .tgt_req(apb_mstr_r1_req),                                                    // o:1
  .tgt_sop(apb_mstr_r1_sop),                                                    // o:1
  .tgt_eop(apb_mstr_r1_eop),                                                    // o:1
  .tgt_flitdata(apb_mstr_r1_flitdata),                                          // o:24
  .tgt_ready(apb_mstr_r1_ready)                                                 // i:1
);
// ============================================================================
// Initiator Port 1 Forward Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Initiator Port 1 Forward Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_f0_dec RTR_INI0_f0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .trigger(trigger),                                                            // i:1
  .ini_activity(RTR_INI0_f0_activity),                                          // i:1
  .ini_req(RTR_INI0_f0_req),                                                    // i:1
  .ini_sop(RTR_INI0_f0_sop),                                                    // i:1
  .ini_eop(RTR_INI0_f0_eop),                                                    // i:1
  .ini_flitdata(RTR_INI0_f0_flitdata),                                          // i:36
  .ini_ready(RTR_INI0_f0_ready),                                                // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // o:1
  .f0_i1_eop(f0_i1_eop),                                                        // o:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // o:4
  .f0_i1_qos(f0_i1_qos),                                                        // o:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // o:36
  .f0_i1_t4_activity(f0_i1_t4_activity),                                        // o:1
  .f0_i1_t4_req_nxt(f0_i1_t4_req_nxt),                                          // o:1
  .f0_i1_t4_req(f0_i1_t4_req),                                                  // o:1
  .f0_i1_t4_ready(f0_i1_t4_ready),                                              // i:1
  .f0_i1_t2_activity(f0_i1_t2_activity),                                        // o:1
  .f0_i1_t2_req_nxt(f0_i1_t2_req_nxt),                                          // o:1
  .f0_i1_t2_req(f0_i1_t2_req),                                                  // o:1
  .f0_i1_t2_ready(f0_i1_t2_ready),                                              // i:1
  .f0_i1_t1_activity(f0_i1_t1_activity),                                        // o:1
  .f0_i1_t1_req_nxt(f0_i1_t1_req_nxt),                                          // o:1
  .f0_i1_t1_req(f0_i1_t1_req),                                                  // o:1
  .f0_i1_t1_ready(f0_i1_t1_ready),                                              // i:1
  .f0_i1_t0_activity(f0_i1_t0_activity),                                        // o:1
  .f0_i1_t0_req_nxt(f0_i1_t0_req_nxt),                                          // o:1
  .f0_i1_t0_req(f0_i1_t0_req),                                                  // o:1
  .f0_i1_t0_ready(f0_i1_t0_ready),                                              // i:1
  .f0_i1_t5_activity(f0_i1_t5_activity),                                        // o:1
  .f0_i1_t5_req_nxt(f0_i1_t5_req_nxt),                                          // o:1
  .f0_i1_t5_req(f0_i1_t5_req),                                                  // o:1
  .f0_i1_t5_ready(f0_i1_t5_ready),                                              // i:1
  .f0_i1_t3_activity(f0_i1_t3_activity),                                        // o:1
  .f0_i1_t3_req_nxt(f0_i1_t3_req_nxt),                                          // o:1
  .f0_i1_t3_req(f0_i1_t3_req),                                                  // o:1
  .f0_i1_t3_ready(f0_i1_t3_ready),                                              // i:1
  .f0_i1_t1000_activity(f0_i1_t1000_activity),                                  // o:1
  .f0_i1_t1000_req_nxt(f0_i1_t1000_req_nxt),                                    // o:1
  .f0_i1_t1000_req(f0_i1_t1000_req),                                            // o:1
  .f0_i1_t1000_ready(f0_i1_t1000_ready)                                         // i:1
);
// ============================================================================
// Initiator Port 1 Forward Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Initiator Port 1 Forward Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_f1_dec RTR_INI0_f1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .trigger(trigger),                                                            // i:1
  .ini_activity(RTR_INI0_f1_activity),                                          // i:1
  .ini_req(RTR_INI0_f1_req),                                                    // i:1
  .ini_sop(RTR_INI0_f1_sop),                                                    // i:1
  .ini_eop(RTR_INI0_f1_eop),                                                    // i:1
  .ini_flitdata(RTR_INI0_f1_flitdata),                                          // i:60
  .ini_ready(RTR_INI0_f1_ready),                                                // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // o:1
  .f1_i1_eop(f1_i1_eop),                                                        // o:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // o:4
  .f1_i1_qos(f1_i1_qos),                                                        // o:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // o:60
  .f1_i1_t4_activity(f1_i1_t4_activity),                                        // o:1
  .f1_i1_t4_req_nxt(f1_i1_t4_req_nxt),                                          // o:1
  .f1_i1_t4_req(f1_i1_t4_req),                                                  // o:1
  .f1_i1_t4_ready(f1_i1_t4_ready),                                              // i:1
  .f1_i1_t2_activity(f1_i1_t2_activity),                                        // o:1
  .f1_i1_t2_req_nxt(f1_i1_t2_req_nxt),                                          // o:1
  .f1_i1_t2_req(f1_i1_t2_req),                                                  // o:1
  .f1_i1_t2_ready(f1_i1_t2_ready),                                              // i:1
  .f1_i1_t1_activity(f1_i1_t1_activity),                                        // o:1
  .f1_i1_t1_req_nxt(f1_i1_t1_req_nxt),                                          // o:1
  .f1_i1_t1_req(f1_i1_t1_req),                                                  // o:1
  .f1_i1_t1_ready(f1_i1_t1_ready),                                              // i:1
  .f1_i1_t0_activity(f1_i1_t0_activity),                                        // o:1
  .f1_i1_t0_req_nxt(f1_i1_t0_req_nxt),                                          // o:1
  .f1_i1_t0_req(f1_i1_t0_req),                                                  // o:1
  .f1_i1_t0_ready(f1_i1_t0_ready),                                              // i:1
  .f1_i1_t5_activity(f1_i1_t5_activity),                                        // o:1
  .f1_i1_t5_req_nxt(f1_i1_t5_req_nxt),                                          // o:1
  .f1_i1_t5_req(f1_i1_t5_req),                                                  // o:1
  .f1_i1_t5_ready(f1_i1_t5_ready),                                              // i:1
  .f1_i1_t3_activity(f1_i1_t3_activity),                                        // o:1
  .f1_i1_t3_req_nxt(f1_i1_t3_req_nxt),                                          // o:1
  .f1_i1_t3_req(f1_i1_t3_req),                                                  // o:1
  .f1_i1_t3_ready(f1_i1_t3_ready),                                              // i:1
  .f1_i1_t1000_activity(f1_i1_t1000_activity),                                  // o:1
  .f1_i1_t1000_req_nxt(f1_i1_t1000_req_nxt),                                    // o:1
  .f1_i1_t1000_req(f1_i1_t1000_req),                                            // o:1
  .f1_i1_t1000_ready(f1_i1_t1000_ready)                                         // i:1
);
// ============================================================================
// Initiator Port 1 Reverse Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Initiator Port 1 Reverse Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_r0_arb RTR_INI0_r0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .r0_t4_sop(r0_t4_sop),                                                        // i:1
  .r0_t4_eop(r0_t4_eop),                                                        // i:1
  .r0_t4_qos_nxt(r0_t4_qos_nxt),                                                // i:4
  .r0_t4_qos(r0_t4_qos),                                                        // i:4
  .r0_t4_flitdata(r0_t4_flitdata),                                              // i:34
  .r0_t4_i1_activity(r0_t4_i1_activity),                                        // i:1
  .r0_t4_i1_req_nxt(r0_t4_i1_req_nxt),                                          // i:1
  .r0_t4_i1_req(r0_t4_i1_req),                                                  // i:1
  .r0_t4_i1_ready(r0_t4_i1_ready),                                              // o:1
  .r0_t2_sop(r0_t2_sop),                                                        // i:1
  .r0_t2_eop(r0_t2_eop),                                                        // i:1
  .r0_t2_qos_nxt(r0_t2_qos_nxt),                                                // i:4
  .r0_t2_qos(r0_t2_qos),                                                        // i:4
  .r0_t2_flitdata(r0_t2_flitdata),                                              // i:34
  .r0_t2_i1_activity(r0_t2_i1_activity),                                        // i:1
  .r0_t2_i1_req_nxt(r0_t2_i1_req_nxt),                                          // i:1
  .r0_t2_i1_req(r0_t2_i1_req),                                                  // i:1
  .r0_t2_i1_ready(r0_t2_i1_ready),                                              // o:1
  .r0_t1_sop(r0_t1_sop),                                                        // i:1
  .r0_t1_eop(r0_t1_eop),                                                        // i:1
  .r0_t1_qos_nxt(r0_t1_qos_nxt),                                                // i:4
  .r0_t1_qos(r0_t1_qos),                                                        // i:4
  .r0_t1_flitdata(r0_t1_flitdata),                                              // i:34
  .r0_t1_i1_activity(r0_t1_i1_activity),                                        // i:1
  .r0_t1_i1_req_nxt(r0_t1_i1_req_nxt),                                          // i:1
  .r0_t1_i1_req(r0_t1_i1_req),                                                  // i:1
  .r0_t1_i1_ready(r0_t1_i1_ready),                                              // o:1
  .r0_t0_sop(r0_t0_sop),                                                        // i:1
  .r0_t0_eop(r0_t0_eop),                                                        // i:1
  .r0_t0_qos_nxt(r0_t0_qos_nxt),                                                // i:4
  .r0_t0_qos(r0_t0_qos),                                                        // i:4
  .r0_t0_flitdata(r0_t0_flitdata),                                              // i:34
  .r0_t0_i1_activity(r0_t0_i1_activity),                                        // i:1
  .r0_t0_i1_req_nxt(r0_t0_i1_req_nxt),                                          // i:1
  .r0_t0_i1_req(r0_t0_i1_req),                                                  // i:1
  .r0_t0_i1_ready(r0_t0_i1_ready),                                              // o:1
  .r0_t5_sop(r0_t5_sop),                                                        // i:1
  .r0_t5_eop(r0_t5_eop),                                                        // i:1
  .r0_t5_qos_nxt(r0_t5_qos_nxt),                                                // i:4
  .r0_t5_qos(r0_t5_qos),                                                        // i:4
  .r0_t5_flitdata(r0_t5_flitdata),                                              // i:34
  .r0_t5_i1_activity(r0_t5_i1_activity),                                        // i:1
  .r0_t5_i1_req_nxt(r0_t5_i1_req_nxt),                                          // i:1
  .r0_t5_i1_req(r0_t5_i1_req),                                                  // i:1
  .r0_t5_i1_ready(r0_t5_i1_ready),                                              // o:1
  .r0_t3_sop(r0_t3_sop),                                                        // i:1
  .r0_t3_eop(r0_t3_eop),                                                        // i:1
  .r0_t3_qos_nxt(r0_t3_qos_nxt),                                                // i:4
  .r0_t3_qos(r0_t3_qos),                                                        // i:4
  .r0_t3_flitdata(r0_t3_flitdata),                                              // i:34
  .r0_t3_i1_activity(r0_t3_i1_activity),                                        // i:1
  .r0_t3_i1_req_nxt(r0_t3_i1_req_nxt),                                          // i:1
  .r0_t3_i1_req(r0_t3_i1_req),                                                  // i:1
  .r0_t3_i1_ready(r0_t3_i1_ready),                                              // o:1
  .r0_t1000_sop(r0_t1000_sop),                                                  // i:1
  .r0_t1000_eop(r0_t1000_eop),                                                  // i:1
  .r0_t1000_qos_nxt(r0_t1000_qos_nxt),                                          // i:4
  .r0_t1000_qos(r0_t1000_qos),                                                  // i:4
  .r0_t1000_flitdata(r0_t1000_flitdata),                                        // i:34
  .r0_t1000_i1_activity(r0_t1000_i1_activity),                                  // i:1
  .r0_t1000_i1_req_nxt(r0_t1000_i1_req_nxt),                                    // i:1
  .r0_t1000_i1_req(r0_t1000_i1_req),                                            // i:1
  .r0_t1000_i1_ready(r0_t1000_i1_ready),                                        // o:1
  .tgt_activity(RTR_INI0_r0_activity),                                          // o:1
  .tgt_req(RTR_INI0_r0_req),                                                    // o:1
  .tgt_sop(RTR_INI0_r0_sop),                                                    // o:1
  .tgt_eop(RTR_INI0_r0_eop),                                                    // o:1
  .tgt_flitdata(RTR_INI0_r0_flitdata),                                          // o:34
  .tgt_ready(RTR_INI0_r0_ready)                                                 // i:1
);
// ============================================================================
// Initiator Port 1 Reverse Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Initiator Port 1 Reverse Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_r1_arb RTR_INI0_r1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .r1_t4_sop(r1_t4_sop),                                                        // i:1
  .r1_t4_eop(r1_t4_eop),                                                        // i:1
  .r1_t4_qos_nxt(r1_t4_qos_nxt),                                                // i:4
  .r1_t4_qos(r1_t4_qos),                                                        // i:4
  .r1_t4_flitdata(r1_t4_flitdata),                                              // i:24
  .r1_t4_i1_activity(r1_t4_i1_activity),                                        // i:1
  .r1_t4_i1_req_nxt(r1_t4_i1_req_nxt),                                          // i:1
  .r1_t4_i1_req(r1_t4_i1_req),                                                  // i:1
  .r1_t4_i1_ready(r1_t4_i1_ready),                                              // o:1
  .r1_t2_sop(r1_t2_sop),                                                        // i:1
  .r1_t2_eop(r1_t2_eop),                                                        // i:1
  .r1_t2_qos_nxt(r1_t2_qos_nxt),                                                // i:4
  .r1_t2_qos(r1_t2_qos),                                                        // i:4
  .r1_t2_flitdata(r1_t2_flitdata),                                              // i:24
  .r1_t2_i1_activity(r1_t2_i1_activity),                                        // i:1
  .r1_t2_i1_req_nxt(r1_t2_i1_req_nxt),                                          // i:1
  .r1_t2_i1_req(r1_t2_i1_req),                                                  // i:1
  .r1_t2_i1_ready(r1_t2_i1_ready),                                              // o:1
  .r1_t1_sop(r1_t1_sop),                                                        // i:1
  .r1_t1_eop(r1_t1_eop),                                                        // i:1
  .r1_t1_qos_nxt(r1_t1_qos_nxt),                                                // i:4
  .r1_t1_qos(r1_t1_qos),                                                        // i:4
  .r1_t1_flitdata(r1_t1_flitdata),                                              // i:24
  .r1_t1_i1_activity(r1_t1_i1_activity),                                        // i:1
  .r1_t1_i1_req_nxt(r1_t1_i1_req_nxt),                                          // i:1
  .r1_t1_i1_req(r1_t1_i1_req),                                                  // i:1
  .r1_t1_i1_ready(r1_t1_i1_ready),                                              // o:1
  .r1_t0_sop(r1_t0_sop),                                                        // i:1
  .r1_t0_eop(r1_t0_eop),                                                        // i:1
  .r1_t0_qos_nxt(r1_t0_qos_nxt),                                                // i:4
  .r1_t0_qos(r1_t0_qos),                                                        // i:4
  .r1_t0_flitdata(r1_t0_flitdata),                                              // i:24
  .r1_t0_i1_activity(r1_t0_i1_activity),                                        // i:1
  .r1_t0_i1_req_nxt(r1_t0_i1_req_nxt),                                          // i:1
  .r1_t0_i1_req(r1_t0_i1_req),                                                  // i:1
  .r1_t0_i1_ready(r1_t0_i1_ready),                                              // o:1
  .r1_t5_sop(r1_t5_sop),                                                        // i:1
  .r1_t5_eop(r1_t5_eop),                                                        // i:1
  .r1_t5_qos_nxt(r1_t5_qos_nxt),                                                // i:4
  .r1_t5_qos(r1_t5_qos),                                                        // i:4
  .r1_t5_flitdata(r1_t5_flitdata),                                              // i:24
  .r1_t5_i1_activity(r1_t5_i1_activity),                                        // i:1
  .r1_t5_i1_req_nxt(r1_t5_i1_req_nxt),                                          // i:1
  .r1_t5_i1_req(r1_t5_i1_req),                                                  // i:1
  .r1_t5_i1_ready(r1_t5_i1_ready),                                              // o:1
  .r1_t3_sop(r1_t3_sop),                                                        // i:1
  .r1_t3_eop(r1_t3_eop),                                                        // i:1
  .r1_t3_qos_nxt(r1_t3_qos_nxt),                                                // i:4
  .r1_t3_qos(r1_t3_qos),                                                        // i:4
  .r1_t3_flitdata(r1_t3_flitdata),                                              // i:24
  .r1_t3_i1_activity(r1_t3_i1_activity),                                        // i:1
  .r1_t3_i1_req_nxt(r1_t3_i1_req_nxt),                                          // i:1
  .r1_t3_i1_req(r1_t3_i1_req),                                                  // i:1
  .r1_t3_i1_ready(r1_t3_i1_ready),                                              // o:1
  .r1_t1000_sop(r1_t1000_sop),                                                  // i:1
  .r1_t1000_eop(r1_t1000_eop),                                                  // i:1
  .r1_t1000_qos_nxt(r1_t1000_qos_nxt),                                          // i:4
  .r1_t1000_qos(r1_t1000_qos),                                                  // i:4
  .r1_t1000_flitdata(r1_t1000_flitdata),                                        // i:24
  .r1_t1000_i1_activity(r1_t1000_i1_activity),                                  // i:1
  .r1_t1000_i1_req_nxt(r1_t1000_i1_req_nxt),                                    // i:1
  .r1_t1000_i1_req(r1_t1000_i1_req),                                            // i:1
  .r1_t1000_i1_ready(r1_t1000_i1_ready),                                        // o:1
  .tgt_activity(RTR_INI0_r1_activity),                                          // o:1
  .tgt_req(RTR_INI0_r1_req),                                                    // o:1
  .tgt_sop(RTR_INI0_r1_sop),                                                    // o:1
  .tgt_eop(RTR_INI0_r1_eop),                                                    // o:1
  .tgt_flitdata(RTR_INI0_r1_flitdata),                                          // o:24
  .tgt_ready(RTR_INI0_r1_ready)                                                 // i:1
);
// ============================================================================
// ============================================================================
// Target Interfaces
// ============================================================================
// ============================================================================
// ============================================================================
// Target Port 0 Forward Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 0 Forward Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb pam3_cmn_TEA_f0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f0_i0_sop(f0_i0_sop),                                                        // i:1
  .f0_i0_eop(f0_i0_eop),                                                        // i:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // i:4
  .f0_i0_qos(f0_i0_qos),                                                        // i:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // i:36
  .f0_i0_t0_activity(f0_i0_t0_activity),                                        // i:1
  .f0_i0_t0_req_nxt(f0_i0_t0_req_nxt),                                          // i:1
  .f0_i0_t0_req(f0_i0_t0_req),                                                  // i:1
  .f0_i0_t0_ready(f0_i0_t0_ready),                                              // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // i:1
  .f0_i1_eop(f0_i1_eop),                                                        // i:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // i:4
  .f0_i1_qos(f0_i1_qos),                                                        // i:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // i:36
  .f0_i1_t0_activity(f0_i1_t0_activity),                                        // i:1
  .f0_i1_t0_req_nxt(f0_i1_t0_req_nxt),                                          // i:1
  .f0_i1_t0_req(f0_i1_t0_req),                                                  // i:1
  .f0_i1_t0_ready(f0_i1_t0_ready),                                              // o:1
  .tgt_activity(pam3_cmn_TEA_f0_activity),                                      // o:1
  .tgt_req(pam3_cmn_TEA_f0_req),                                                // o:1
  .tgt_sop(pam3_cmn_TEA_f0_sop),                                                // o:1
  .tgt_eop(pam3_cmn_TEA_f0_eop),                                                // o:1
  .tgt_flitdata(pam3_cmn_TEA_f0_flitdata),                                      // o:36
  .tgt_ready(pam3_cmn_TEA_f0_ready)                                             // i:1
);
// ============================================================================
// Target Port 0 Forward Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 0 Forward Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb pam3_cmn_TEA_f1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f1_i0_sop(f1_i0_sop),                                                        // i:1
  .f1_i0_eop(f1_i0_eop),                                                        // i:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // i:4
  .f1_i0_qos(f1_i0_qos),                                                        // i:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // i:60
  .f1_i0_t0_activity(f1_i0_t0_activity),                                        // i:1
  .f1_i0_t0_req_nxt(f1_i0_t0_req_nxt),                                          // i:1
  .f1_i0_t0_req(f1_i0_t0_req),                                                  // i:1
  .f1_i0_t0_ready(f1_i0_t0_ready),                                              // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // i:1
  .f1_i1_eop(f1_i1_eop),                                                        // i:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // i:4
  .f1_i1_qos(f1_i1_qos),                                                        // i:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // i:60
  .f1_i1_t0_activity(f1_i1_t0_activity),                                        // i:1
  .f1_i1_t0_req_nxt(f1_i1_t0_req_nxt),                                          // i:1
  .f1_i1_t0_req(f1_i1_t0_req),                                                  // i:1
  .f1_i1_t0_ready(f1_i1_t0_ready),                                              // o:1
  .tgt_activity(pam3_cmn_TEA_f1_activity),                                      // o:1
  .tgt_req(pam3_cmn_TEA_f1_req),                                                // o:1
  .tgt_sop(pam3_cmn_TEA_f1_sop),                                                // o:1
  .tgt_eop(pam3_cmn_TEA_f1_eop),                                                // o:1
  .tgt_flitdata(pam3_cmn_TEA_f1_flitdata),                                      // o:60
  .tgt_ready(pam3_cmn_TEA_f1_ready)                                             // i:1
);
// ============================================================================
// Target Port 0 Reverse Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 0 Reverse Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec pam3_cmn_TEA_r0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(pam3_cmn_TEA_r0_activity),                                      // i:1
  .ini_req(pam3_cmn_TEA_r0_req),                                                // i:1
  .ini_sop(pam3_cmn_TEA_r0_sop),                                                // i:1
  .ini_eop(pam3_cmn_TEA_r0_eop),                                                // i:1
  .ini_flitdata(pam3_cmn_TEA_r0_flitdata),                                      // i:34
  .ini_ready(pam3_cmn_TEA_r0_ready),                                            // o:1
  .r0_t0_sop(r0_t0_sop),                                                        // o:1
  .r0_t0_eop(r0_t0_eop),                                                        // o:1
  .r0_t0_qos_nxt(r0_t0_qos_nxt),                                                // o:4
  .r0_t0_qos(r0_t0_qos),                                                        // o:4
  .r0_t0_flitdata(r0_t0_flitdata),                                              // o:34
  .r0_t0_i0_activity(r0_t0_i0_activity),                                        // o:1
  .r0_t0_i0_req_nxt(r0_t0_i0_req_nxt),                                          // o:1
  .r0_t0_i0_req(r0_t0_i0_req),                                                  // o:1
  .r0_t0_i0_ready(r0_t0_i0_ready),                                              // i:1
  .r0_t0_i1_activity(r0_t0_i1_activity),                                        // o:1
  .r0_t0_i1_req_nxt(r0_t0_i1_req_nxt),                                          // o:1
  .r0_t0_i1_req(r0_t0_i1_req),                                                  // o:1
  .r0_t0_i1_ready(r0_t0_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 0 Reverse Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 0 Reverse Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec pam3_cmn_TEA_r1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(pam3_cmn_TEA_r1_activity),                                      // i:1
  .ini_req(pam3_cmn_TEA_r1_req),                                                // i:1
  .ini_sop(pam3_cmn_TEA_r1_sop),                                                // i:1
  .ini_eop(pam3_cmn_TEA_r1_eop),                                                // i:1
  .ini_flitdata(pam3_cmn_TEA_r1_flitdata),                                      // i:24
  .ini_ready(pam3_cmn_TEA_r1_ready),                                            // o:1
  .r1_t0_sop(r1_t0_sop),                                                        // o:1
  .r1_t0_eop(r1_t0_eop),                                                        // o:1
  .r1_t0_qos_nxt(r1_t0_qos_nxt),                                                // o:4
  .r1_t0_qos(r1_t0_qos),                                                        // o:4
  .r1_t0_flitdata(r1_t0_flitdata),                                              // o:24
  .r1_t0_i0_activity(r1_t0_i0_activity),                                        // o:1
  .r1_t0_i0_req_nxt(r1_t0_i0_req_nxt),                                          // o:1
  .r1_t0_i0_req(r1_t0_i0_req),                                                  // o:1
  .r1_t0_i0_ready(r1_t0_i0_ready),                                              // i:1
  .r1_t0_i1_activity(r1_t0_i1_activity),                                        // o:1
  .r1_t0_i1_req_nxt(r1_t0_i1_req_nxt),                                          // o:1
  .r1_t0_i1_req(r1_t0_i1_req),                                                  // o:1
  .r1_t0_i1_ready(r1_t0_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 1 Forward Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 1 Forward Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb tc_reg_TEA_f0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f0_i0_sop(f0_i0_sop),                                                        // i:1
  .f0_i0_eop(f0_i0_eop),                                                        // i:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // i:4
  .f0_i0_qos(f0_i0_qos),                                                        // i:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // i:36
  .f0_i0_t1_activity(f0_i0_t1_activity),                                        // i:1
  .f0_i0_t1_req_nxt(f0_i0_t1_req_nxt),                                          // i:1
  .f0_i0_t1_req(f0_i0_t1_req),                                                  // i:1
  .f0_i0_t1_ready(f0_i0_t1_ready),                                              // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // i:1
  .f0_i1_eop(f0_i1_eop),                                                        // i:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // i:4
  .f0_i1_qos(f0_i1_qos),                                                        // i:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // i:36
  .f0_i1_t1_activity(f0_i1_t1_activity),                                        // i:1
  .f0_i1_t1_req_nxt(f0_i1_t1_req_nxt),                                          // i:1
  .f0_i1_t1_req(f0_i1_t1_req),                                                  // i:1
  .f0_i1_t1_ready(f0_i1_t1_ready),                                              // o:1
  .tgt_activity(tc_reg_TEA_f0_activity),                                        // o:1
  .tgt_req(tc_reg_TEA_f0_req),                                                  // o:1
  .tgt_sop(tc_reg_TEA_f0_sop),                                                  // o:1
  .tgt_eop(tc_reg_TEA_f0_eop),                                                  // o:1
  .tgt_flitdata(tc_reg_TEA_f0_flitdata),                                        // o:36
  .tgt_ready(tc_reg_TEA_f0_ready)                                               // i:1
);
// ============================================================================
// Target Port 1 Forward Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 1 Forward Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb tc_reg_TEA_f1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f1_i0_sop(f1_i0_sop),                                                        // i:1
  .f1_i0_eop(f1_i0_eop),                                                        // i:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // i:4
  .f1_i0_qos(f1_i0_qos),                                                        // i:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // i:60
  .f1_i0_t1_activity(f1_i0_t1_activity),                                        // i:1
  .f1_i0_t1_req_nxt(f1_i0_t1_req_nxt),                                          // i:1
  .f1_i0_t1_req(f1_i0_t1_req),                                                  // i:1
  .f1_i0_t1_ready(f1_i0_t1_ready),                                              // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // i:1
  .f1_i1_eop(f1_i1_eop),                                                        // i:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // i:4
  .f1_i1_qos(f1_i1_qos),                                                        // i:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // i:60
  .f1_i1_t1_activity(f1_i1_t1_activity),                                        // i:1
  .f1_i1_t1_req_nxt(f1_i1_t1_req_nxt),                                          // i:1
  .f1_i1_t1_req(f1_i1_t1_req),                                                  // i:1
  .f1_i1_t1_ready(f1_i1_t1_ready),                                              // o:1
  .tgt_activity(tc_reg_TEA_f1_activity),                                        // o:1
  .tgt_req(tc_reg_TEA_f1_req),                                                  // o:1
  .tgt_sop(tc_reg_TEA_f1_sop),                                                  // o:1
  .tgt_eop(tc_reg_TEA_f1_eop),                                                  // o:1
  .tgt_flitdata(tc_reg_TEA_f1_flitdata),                                        // o:60
  .tgt_ready(tc_reg_TEA_f1_ready)                                               // i:1
);
// ============================================================================
// Target Port 1 Reverse Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 1 Reverse Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec tc_reg_TEA_r0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(tc_reg_TEA_r0_activity),                                        // i:1
  .ini_req(tc_reg_TEA_r0_req),                                                  // i:1
  .ini_sop(tc_reg_TEA_r0_sop),                                                  // i:1
  .ini_eop(tc_reg_TEA_r0_eop),                                                  // i:1
  .ini_flitdata(tc_reg_TEA_r0_flitdata),                                        // i:34
  .ini_ready(tc_reg_TEA_r0_ready),                                              // o:1
  .r0_t1_sop(r0_t1_sop),                                                        // o:1
  .r0_t1_eop(r0_t1_eop),                                                        // o:1
  .r0_t1_qos_nxt(r0_t1_qos_nxt),                                                // o:4
  .r0_t1_qos(r0_t1_qos),                                                        // o:4
  .r0_t1_flitdata(r0_t1_flitdata),                                              // o:34
  .r0_t1_i0_activity(r0_t1_i0_activity),                                        // o:1
  .r0_t1_i0_req_nxt(r0_t1_i0_req_nxt),                                          // o:1
  .r0_t1_i0_req(r0_t1_i0_req),                                                  // o:1
  .r0_t1_i0_ready(r0_t1_i0_ready),                                              // i:1
  .r0_t1_i1_activity(r0_t1_i1_activity),                                        // o:1
  .r0_t1_i1_req_nxt(r0_t1_i1_req_nxt),                                          // o:1
  .r0_t1_i1_req(r0_t1_i1_req),                                                  // o:1
  .r0_t1_i1_ready(r0_t1_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 1 Reverse Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 1 Reverse Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec tc_reg_TEA_r1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(tc_reg_TEA_r1_activity),                                        // i:1
  .ini_req(tc_reg_TEA_r1_req),                                                  // i:1
  .ini_sop(tc_reg_TEA_r1_sop),                                                  // i:1
  .ini_eop(tc_reg_TEA_r1_eop),                                                  // i:1
  .ini_flitdata(tc_reg_TEA_r1_flitdata),                                        // i:24
  .ini_ready(tc_reg_TEA_r1_ready),                                              // o:1
  .r1_t1_sop(r1_t1_sop),                                                        // o:1
  .r1_t1_eop(r1_t1_eop),                                                        // o:1
  .r1_t1_qos_nxt(r1_t1_qos_nxt),                                                // o:4
  .r1_t1_qos(r1_t1_qos),                                                        // o:4
  .r1_t1_flitdata(r1_t1_flitdata),                                              // o:24
  .r1_t1_i0_activity(r1_t1_i0_activity),                                        // o:1
  .r1_t1_i0_req_nxt(r1_t1_i0_req_nxt),                                          // o:1
  .r1_t1_i0_req(r1_t1_i0_req),                                                  // o:1
  .r1_t1_i0_ready(r1_t1_i0_ready),                                              // i:1
  .r1_t1_i1_activity(r1_t1_i1_activity),                                        // o:1
  .r1_t1_i1_req_nxt(r1_t1_i1_req_nxt),                                          // o:1
  .r1_t1_i1_req(r1_t1_i1_req),                                                  // o:1
  .r1_t1_i1_ready(r1_t1_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 2 Forward Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 2 Forward Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb usb_sub_sys_TEA_f0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f0_i0_sop(f0_i0_sop),                                                        // i:1
  .f0_i0_eop(f0_i0_eop),                                                        // i:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // i:4
  .f0_i0_qos(f0_i0_qos),                                                        // i:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // i:36
  .f0_i0_t2_activity(f0_i0_t2_activity),                                        // i:1
  .f0_i0_t2_req_nxt(f0_i0_t2_req_nxt),                                          // i:1
  .f0_i0_t2_req(f0_i0_t2_req),                                                  // i:1
  .f0_i0_t2_ready(f0_i0_t2_ready),                                              // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // i:1
  .f0_i1_eop(f0_i1_eop),                                                        // i:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // i:4
  .f0_i1_qos(f0_i1_qos),                                                        // i:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // i:36
  .f0_i1_t2_activity(f0_i1_t2_activity),                                        // i:1
  .f0_i1_t2_req_nxt(f0_i1_t2_req_nxt),                                          // i:1
  .f0_i1_t2_req(f0_i1_t2_req),                                                  // i:1
  .f0_i1_t2_ready(f0_i1_t2_ready),                                              // o:1
  .tgt_activity(usb_sub_sys_TEA_f0_activity),                                   // o:1
  .tgt_req(usb_sub_sys_TEA_f0_req),                                             // o:1
  .tgt_sop(usb_sub_sys_TEA_f0_sop),                                             // o:1
  .tgt_eop(usb_sub_sys_TEA_f0_eop),                                             // o:1
  .tgt_flitdata(usb_sub_sys_TEA_f0_flitdata),                                   // o:36
  .tgt_ready(usb_sub_sys_TEA_f0_ready)                                          // i:1
);
// ============================================================================
// Target Port 2 Forward Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 2 Forward Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb usb_sub_sys_TEA_f1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f1_i0_sop(f1_i0_sop),                                                        // i:1
  .f1_i0_eop(f1_i0_eop),                                                        // i:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // i:4
  .f1_i0_qos(f1_i0_qos),                                                        // i:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // i:60
  .f1_i0_t2_activity(f1_i0_t2_activity),                                        // i:1
  .f1_i0_t2_req_nxt(f1_i0_t2_req_nxt),                                          // i:1
  .f1_i0_t2_req(f1_i0_t2_req),                                                  // i:1
  .f1_i0_t2_ready(f1_i0_t2_ready),                                              // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // i:1
  .f1_i1_eop(f1_i1_eop),                                                        // i:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // i:4
  .f1_i1_qos(f1_i1_qos),                                                        // i:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // i:60
  .f1_i1_t2_activity(f1_i1_t2_activity),                                        // i:1
  .f1_i1_t2_req_nxt(f1_i1_t2_req_nxt),                                          // i:1
  .f1_i1_t2_req(f1_i1_t2_req),                                                  // i:1
  .f1_i1_t2_ready(f1_i1_t2_ready),                                              // o:1
  .tgt_activity(usb_sub_sys_TEA_f1_activity),                                   // o:1
  .tgt_req(usb_sub_sys_TEA_f1_req),                                             // o:1
  .tgt_sop(usb_sub_sys_TEA_f1_sop),                                             // o:1
  .tgt_eop(usb_sub_sys_TEA_f1_eop),                                             // o:1
  .tgt_flitdata(usb_sub_sys_TEA_f1_flitdata),                                   // o:60
  .tgt_ready(usb_sub_sys_TEA_f1_ready)                                          // i:1
);
// ============================================================================
// Target Port 2 Reverse Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 2 Reverse Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec usb_sub_sys_TEA_r0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(usb_sub_sys_TEA_r0_activity),                                   // i:1
  .ini_req(usb_sub_sys_TEA_r0_req),                                             // i:1
  .ini_sop(usb_sub_sys_TEA_r0_sop),                                             // i:1
  .ini_eop(usb_sub_sys_TEA_r0_eop),                                             // i:1
  .ini_flitdata(usb_sub_sys_TEA_r0_flitdata),                                   // i:34
  .ini_ready(usb_sub_sys_TEA_r0_ready),                                         // o:1
  .r0_t2_sop(r0_t2_sop),                                                        // o:1
  .r0_t2_eop(r0_t2_eop),                                                        // o:1
  .r0_t2_qos_nxt(r0_t2_qos_nxt),                                                // o:4
  .r0_t2_qos(r0_t2_qos),                                                        // o:4
  .r0_t2_flitdata(r0_t2_flitdata),                                              // o:34
  .r0_t2_i0_activity(r0_t2_i0_activity),                                        // o:1
  .r0_t2_i0_req_nxt(r0_t2_i0_req_nxt),                                          // o:1
  .r0_t2_i0_req(r0_t2_i0_req),                                                  // o:1
  .r0_t2_i0_ready(r0_t2_i0_ready),                                              // i:1
  .r0_t2_i1_activity(r0_t2_i1_activity),                                        // o:1
  .r0_t2_i1_req_nxt(r0_t2_i1_req_nxt),                                          // o:1
  .r0_t2_i1_req(r0_t2_i1_req),                                                  // o:1
  .r0_t2_i1_ready(r0_t2_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 2 Reverse Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 2 Reverse Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec usb_sub_sys_TEA_r1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(usb_sub_sys_TEA_r1_activity),                                   // i:1
  .ini_req(usb_sub_sys_TEA_r1_req),                                             // i:1
  .ini_sop(usb_sub_sys_TEA_r1_sop),                                             // i:1
  .ini_eop(usb_sub_sys_TEA_r1_eop),                                             // i:1
  .ini_flitdata(usb_sub_sys_TEA_r1_flitdata),                                   // i:24
  .ini_ready(usb_sub_sys_TEA_r1_ready),                                         // o:1
  .r1_t2_sop(r1_t2_sop),                                                        // o:1
  .r1_t2_eop(r1_t2_eop),                                                        // o:1
  .r1_t2_qos_nxt(r1_t2_qos_nxt),                                                // o:4
  .r1_t2_qos(r1_t2_qos),                                                        // o:4
  .r1_t2_flitdata(r1_t2_flitdata),                                              // o:24
  .r1_t2_i0_activity(r1_t2_i0_activity),                                        // o:1
  .r1_t2_i0_req_nxt(r1_t2_i0_req_nxt),                                          // o:1
  .r1_t2_i0_req(r1_t2_i0_req),                                                  // o:1
  .r1_t2_i0_ready(r1_t2_i0_ready),                                              // i:1
  .r1_t2_i1_activity(r1_t2_i1_activity),                                        // o:1
  .r1_t2_i1_req_nxt(r1_t2_i1_req_nxt),                                          // o:1
  .r1_t2_i1_req(r1_t2_i1_req),                                                  // o:1
  .r1_t2_i1_ready(r1_t2_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 3 Forward Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 3 Forward Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb pam3_sub_sys_TEA_f0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f0_i0_sop(f0_i0_sop),                                                        // i:1
  .f0_i0_eop(f0_i0_eop),                                                        // i:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // i:4
  .f0_i0_qos(f0_i0_qos),                                                        // i:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // i:36
  .f0_i0_t3_activity(f0_i0_t3_activity),                                        // i:1
  .f0_i0_t3_req_nxt(f0_i0_t3_req_nxt),                                          // i:1
  .f0_i0_t3_req(f0_i0_t3_req),                                                  // i:1
  .f0_i0_t3_ready(f0_i0_t3_ready),                                              // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // i:1
  .f0_i1_eop(f0_i1_eop),                                                        // i:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // i:4
  .f0_i1_qos(f0_i1_qos),                                                        // i:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // i:36
  .f0_i1_t3_activity(f0_i1_t3_activity),                                        // i:1
  .f0_i1_t3_req_nxt(f0_i1_t3_req_nxt),                                          // i:1
  .f0_i1_t3_req(f0_i1_t3_req),                                                  // i:1
  .f0_i1_t3_ready(f0_i1_t3_ready),                                              // o:1
  .tgt_activity(pam3_sub_sys_TEA_f0_activity),                                  // o:1
  .tgt_req(pam3_sub_sys_TEA_f0_req),                                            // o:1
  .tgt_sop(pam3_sub_sys_TEA_f0_sop),                                            // o:1
  .tgt_eop(pam3_sub_sys_TEA_f0_eop),                                            // o:1
  .tgt_flitdata(pam3_sub_sys_TEA_f0_flitdata),                                  // o:36
  .tgt_ready(pam3_sub_sys_TEA_f0_ready)                                         // i:1
);
// ============================================================================
// Target Port 3 Forward Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 3 Forward Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb pam3_sub_sys_TEA_f1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f1_i0_sop(f1_i0_sop),                                                        // i:1
  .f1_i0_eop(f1_i0_eop),                                                        // i:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // i:4
  .f1_i0_qos(f1_i0_qos),                                                        // i:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // i:60
  .f1_i0_t3_activity(f1_i0_t3_activity),                                        // i:1
  .f1_i0_t3_req_nxt(f1_i0_t3_req_nxt),                                          // i:1
  .f1_i0_t3_req(f1_i0_t3_req),                                                  // i:1
  .f1_i0_t3_ready(f1_i0_t3_ready),                                              // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // i:1
  .f1_i1_eop(f1_i1_eop),                                                        // i:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // i:4
  .f1_i1_qos(f1_i1_qos),                                                        // i:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // i:60
  .f1_i1_t3_activity(f1_i1_t3_activity),                                        // i:1
  .f1_i1_t3_req_nxt(f1_i1_t3_req_nxt),                                          // i:1
  .f1_i1_t3_req(f1_i1_t3_req),                                                  // i:1
  .f1_i1_t3_ready(f1_i1_t3_ready),                                              // o:1
  .tgt_activity(pam3_sub_sys_TEA_f1_activity),                                  // o:1
  .tgt_req(pam3_sub_sys_TEA_f1_req),                                            // o:1
  .tgt_sop(pam3_sub_sys_TEA_f1_sop),                                            // o:1
  .tgt_eop(pam3_sub_sys_TEA_f1_eop),                                            // o:1
  .tgt_flitdata(pam3_sub_sys_TEA_f1_flitdata),                                  // o:60
  .tgt_ready(pam3_sub_sys_TEA_f1_ready)                                         // i:1
);
// ============================================================================
// Target Port 3 Reverse Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 3 Reverse Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec pam3_sub_sys_TEA_r0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(pam3_sub_sys_TEA_r0_activity),                                  // i:1
  .ini_req(pam3_sub_sys_TEA_r0_req),                                            // i:1
  .ini_sop(pam3_sub_sys_TEA_r0_sop),                                            // i:1
  .ini_eop(pam3_sub_sys_TEA_r0_eop),                                            // i:1
  .ini_flitdata(pam3_sub_sys_TEA_r0_flitdata),                                  // i:34
  .ini_ready(pam3_sub_sys_TEA_r0_ready),                                        // o:1
  .r0_t3_sop(r0_t3_sop),                                                        // o:1
  .r0_t3_eop(r0_t3_eop),                                                        // o:1
  .r0_t3_qos_nxt(r0_t3_qos_nxt),                                                // o:4
  .r0_t3_qos(r0_t3_qos),                                                        // o:4
  .r0_t3_flitdata(r0_t3_flitdata),                                              // o:34
  .r0_t3_i0_activity(r0_t3_i0_activity),                                        // o:1
  .r0_t3_i0_req_nxt(r0_t3_i0_req_nxt),                                          // o:1
  .r0_t3_i0_req(r0_t3_i0_req),                                                  // o:1
  .r0_t3_i0_ready(r0_t3_i0_ready),                                              // i:1
  .r0_t3_i1_activity(r0_t3_i1_activity),                                        // o:1
  .r0_t3_i1_req_nxt(r0_t3_i1_req_nxt),                                          // o:1
  .r0_t3_i1_req(r0_t3_i1_req),                                                  // o:1
  .r0_t3_i1_ready(r0_t3_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 3 Reverse Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 3 Reverse Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec pam3_sub_sys_TEA_r1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(pam3_sub_sys_TEA_r1_activity),                                  // i:1
  .ini_req(pam3_sub_sys_TEA_r1_req),                                            // i:1
  .ini_sop(pam3_sub_sys_TEA_r1_sop),                                            // i:1
  .ini_eop(pam3_sub_sys_TEA_r1_eop),                                            // i:1
  .ini_flitdata(pam3_sub_sys_TEA_r1_flitdata),                                  // i:24
  .ini_ready(pam3_sub_sys_TEA_r1_ready),                                        // o:1
  .r1_t3_sop(r1_t3_sop),                                                        // o:1
  .r1_t3_eop(r1_t3_eop),                                                        // o:1
  .r1_t3_qos_nxt(r1_t3_qos_nxt),                                                // o:4
  .r1_t3_qos(r1_t3_qos),                                                        // o:4
  .r1_t3_flitdata(r1_t3_flitdata),                                              // o:24
  .r1_t3_i0_activity(r1_t3_i0_activity),                                        // o:1
  .r1_t3_i0_req_nxt(r1_t3_i0_req_nxt),                                          // o:1
  .r1_t3_i0_req(r1_t3_i0_req),                                                  // o:1
  .r1_t3_i0_ready(r1_t3_i0_ready),                                              // i:1
  .r1_t3_i1_activity(r1_t3_i1_activity),                                        // o:1
  .r1_t3_i1_req_nxt(r1_t3_i1_req_nxt),                                          // o:1
  .r1_t3_i1_req(r1_t3_i1_req),                                                  // o:1
  .r1_t3_i1_ready(r1_t3_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 4 Forward Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 4 Forward Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb usb4_phy_TEA_f0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f0_i0_sop(f0_i0_sop),                                                        // i:1
  .f0_i0_eop(f0_i0_eop),                                                        // i:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // i:4
  .f0_i0_qos(f0_i0_qos),                                                        // i:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // i:36
  .f0_i0_t4_activity(f0_i0_t4_activity),                                        // i:1
  .f0_i0_t4_req_nxt(f0_i0_t4_req_nxt),                                          // i:1
  .f0_i0_t4_req(f0_i0_t4_req),                                                  // i:1
  .f0_i0_t4_ready(f0_i0_t4_ready),                                              // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // i:1
  .f0_i1_eop(f0_i1_eop),                                                        // i:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // i:4
  .f0_i1_qos(f0_i1_qos),                                                        // i:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // i:36
  .f0_i1_t4_activity(f0_i1_t4_activity),                                        // i:1
  .f0_i1_t4_req_nxt(f0_i1_t4_req_nxt),                                          // i:1
  .f0_i1_t4_req(f0_i1_t4_req),                                                  // i:1
  .f0_i1_t4_ready(f0_i1_t4_ready),                                              // o:1
  .tgt_activity(usb4_phy_TEA_f0_activity),                                      // o:1
  .tgt_req(usb4_phy_TEA_f0_req),                                                // o:1
  .tgt_sop(usb4_phy_TEA_f0_sop),                                                // o:1
  .tgt_eop(usb4_phy_TEA_f0_eop),                                                // o:1
  .tgt_flitdata(usb4_phy_TEA_f0_flitdata),                                      // o:36
  .tgt_ready(usb4_phy_TEA_f0_ready)                                             // i:1
);
// ============================================================================
// Target Port 4 Forward Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 4 Forward Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb usb4_phy_TEA_f1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f1_i0_sop(f1_i0_sop),                                                        // i:1
  .f1_i0_eop(f1_i0_eop),                                                        // i:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // i:4
  .f1_i0_qos(f1_i0_qos),                                                        // i:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // i:60
  .f1_i0_t4_activity(f1_i0_t4_activity),                                        // i:1
  .f1_i0_t4_req_nxt(f1_i0_t4_req_nxt),                                          // i:1
  .f1_i0_t4_req(f1_i0_t4_req),                                                  // i:1
  .f1_i0_t4_ready(f1_i0_t4_ready),                                              // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // i:1
  .f1_i1_eop(f1_i1_eop),                                                        // i:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // i:4
  .f1_i1_qos(f1_i1_qos),                                                        // i:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // i:60
  .f1_i1_t4_activity(f1_i1_t4_activity),                                        // i:1
  .f1_i1_t4_req_nxt(f1_i1_t4_req_nxt),                                          // i:1
  .f1_i1_t4_req(f1_i1_t4_req),                                                  // i:1
  .f1_i1_t4_ready(f1_i1_t4_ready),                                              // o:1
  .tgt_activity(usb4_phy_TEA_f1_activity),                                      // o:1
  .tgt_req(usb4_phy_TEA_f1_req),                                                // o:1
  .tgt_sop(usb4_phy_TEA_f1_sop),                                                // o:1
  .tgt_eop(usb4_phy_TEA_f1_eop),                                                // o:1
  .tgt_flitdata(usb4_phy_TEA_f1_flitdata),                                      // o:60
  .tgt_ready(usb4_phy_TEA_f1_ready)                                             // i:1
);
// ============================================================================
// Target Port 4 Reverse Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 4 Reverse Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec usb4_phy_TEA_r0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(usb4_phy_TEA_r0_activity),                                      // i:1
  .ini_req(usb4_phy_TEA_r0_req),                                                // i:1
  .ini_sop(usb4_phy_TEA_r0_sop),                                                // i:1
  .ini_eop(usb4_phy_TEA_r0_eop),                                                // i:1
  .ini_flitdata(usb4_phy_TEA_r0_flitdata),                                      // i:34
  .ini_ready(usb4_phy_TEA_r0_ready),                                            // o:1
  .r0_t4_sop(r0_t4_sop),                                                        // o:1
  .r0_t4_eop(r0_t4_eop),                                                        // o:1
  .r0_t4_qos_nxt(r0_t4_qos_nxt),                                                // o:4
  .r0_t4_qos(r0_t4_qos),                                                        // o:4
  .r0_t4_flitdata(r0_t4_flitdata),                                              // o:34
  .r0_t4_i0_activity(r0_t4_i0_activity),                                        // o:1
  .r0_t4_i0_req_nxt(r0_t4_i0_req_nxt),                                          // o:1
  .r0_t4_i0_req(r0_t4_i0_req),                                                  // o:1
  .r0_t4_i0_ready(r0_t4_i0_ready),                                              // i:1
  .r0_t4_i1_activity(r0_t4_i1_activity),                                        // o:1
  .r0_t4_i1_req_nxt(r0_t4_i1_req_nxt),                                          // o:1
  .r0_t4_i1_req(r0_t4_i1_req),                                                  // o:1
  .r0_t4_i1_ready(r0_t4_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 4 Reverse Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 4 Reverse Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec usb4_phy_TEA_r1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(usb4_phy_TEA_r1_activity),                                      // i:1
  .ini_req(usb4_phy_TEA_r1_req),                                                // i:1
  .ini_sop(usb4_phy_TEA_r1_sop),                                                // i:1
  .ini_eop(usb4_phy_TEA_r1_eop),                                                // i:1
  .ini_flitdata(usb4_phy_TEA_r1_flitdata),                                      // i:24
  .ini_ready(usb4_phy_TEA_r1_ready),                                            // o:1
  .r1_t4_sop(r1_t4_sop),                                                        // o:1
  .r1_t4_eop(r1_t4_eop),                                                        // o:1
  .r1_t4_qos_nxt(r1_t4_qos_nxt),                                                // o:4
  .r1_t4_qos(r1_t4_qos),                                                        // o:4
  .r1_t4_flitdata(r1_t4_flitdata),                                              // o:24
  .r1_t4_i0_activity(r1_t4_i0_activity),                                        // o:1
  .r1_t4_i0_req_nxt(r1_t4_i0_req_nxt),                                          // o:1
  .r1_t4_i0_req(r1_t4_i0_req),                                                  // o:1
  .r1_t4_i0_ready(r1_t4_i0_ready),                                              // i:1
  .r1_t4_i1_activity(r1_t4_i1_activity),                                        // o:1
  .r1_t4_i1_req_nxt(r1_t4_i1_req_nxt),                                          // o:1
  .r1_t4_i1_req(r1_t4_i1_req),                                                  // o:1
  .r1_t4_i1_ready(r1_t4_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 5 Forward Channel 0 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 5 Forward Channel 0 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb pam3_xcvr_TEA_f0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f0_i0_sop(f0_i0_sop),                                                        // i:1
  .f0_i0_eop(f0_i0_eop),                                                        // i:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // i:4
  .f0_i0_qos(f0_i0_qos),                                                        // i:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // i:36
  .f0_i0_t5_activity(f0_i0_t5_activity),                                        // i:1
  .f0_i0_t5_req_nxt(f0_i0_t5_req_nxt),                                          // i:1
  .f0_i0_t5_req(f0_i0_t5_req),                                                  // i:1
  .f0_i0_t5_ready(f0_i0_t5_ready),                                              // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // i:1
  .f0_i1_eop(f0_i1_eop),                                                        // i:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // i:4
  .f0_i1_qos(f0_i1_qos),                                                        // i:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // i:36
  .f0_i1_t5_activity(f0_i1_t5_activity),                                        // i:1
  .f0_i1_t5_req_nxt(f0_i1_t5_req_nxt),                                          // i:1
  .f0_i1_t5_req(f0_i1_t5_req),                                                  // i:1
  .f0_i1_t5_ready(f0_i1_t5_ready),                                              // o:1
  .tgt_activity(pam3_xcvr_TEA_f0_activity),                                     // o:1
  .tgt_req(pam3_xcvr_TEA_f0_req),                                               // o:1
  .tgt_sop(pam3_xcvr_TEA_f0_sop),                                               // o:1
  .tgt_eop(pam3_xcvr_TEA_f0_eop),                                               // o:1
  .tgt_flitdata(pam3_xcvr_TEA_f0_flitdata),                                     // o:36
  .tgt_ready(pam3_xcvr_TEA_f0_ready)                                            // i:1
);
// ============================================================================
// Target Port 5 Forward Channel 1 Interface (LLK manager)
// ============================================================================
// ============================================================================
// Target Port 5 Forward Channel 1 Arbiter
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb pam3_xcvr_TEA_f1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .f1_i0_sop(f1_i0_sop),                                                        // i:1
  .f1_i0_eop(f1_i0_eop),                                                        // i:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // i:4
  .f1_i0_qos(f1_i0_qos),                                                        // i:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // i:60
  .f1_i0_t5_activity(f1_i0_t5_activity),                                        // i:1
  .f1_i0_t5_req_nxt(f1_i0_t5_req_nxt),                                          // i:1
  .f1_i0_t5_req(f1_i0_t5_req),                                                  // i:1
  .f1_i0_t5_ready(f1_i0_t5_ready),                                              // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // i:1
  .f1_i1_eop(f1_i1_eop),                                                        // i:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // i:4
  .f1_i1_qos(f1_i1_qos),                                                        // i:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // i:60
  .f1_i1_t5_activity(f1_i1_t5_activity),                                        // i:1
  .f1_i1_t5_req_nxt(f1_i1_t5_req_nxt),                                          // i:1
  .f1_i1_t5_req(f1_i1_t5_req),                                                  // i:1
  .f1_i1_t5_ready(f1_i1_t5_ready),                                              // o:1
  .tgt_activity(pam3_xcvr_TEA_f1_activity),                                     // o:1
  .tgt_req(pam3_xcvr_TEA_f1_req),                                               // o:1
  .tgt_sop(pam3_xcvr_TEA_f1_sop),                                               // o:1
  .tgt_eop(pam3_xcvr_TEA_f1_eop),                                               // o:1
  .tgt_flitdata(pam3_xcvr_TEA_f1_flitdata),                                     // o:60
  .tgt_ready(pam3_xcvr_TEA_f1_ready)                                            // i:1
);
// ============================================================================
// Target Port 5 Reverse Channel 0 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 5 Reverse Channel 0 Decoder
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec pam3_xcvr_TEA_r0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(pam3_xcvr_TEA_r0_activity),                                     // i:1
  .ini_req(pam3_xcvr_TEA_r0_req),                                               // i:1
  .ini_sop(pam3_xcvr_TEA_r0_sop),                                               // i:1
  .ini_eop(pam3_xcvr_TEA_r0_eop),                                               // i:1
  .ini_flitdata(pam3_xcvr_TEA_r0_flitdata),                                     // i:34
  .ini_ready(pam3_xcvr_TEA_r0_ready),                                           // o:1
  .r0_t5_sop(r0_t5_sop),                                                        // o:1
  .r0_t5_eop(r0_t5_eop),                                                        // o:1
  .r0_t5_qos_nxt(r0_t5_qos_nxt),                                                // o:4
  .r0_t5_qos(r0_t5_qos),                                                        // o:4
  .r0_t5_flitdata(r0_t5_flitdata),                                              // o:34
  .r0_t5_i0_activity(r0_t5_i0_activity),                                        // o:1
  .r0_t5_i0_req_nxt(r0_t5_i0_req_nxt),                                          // o:1
  .r0_t5_i0_req(r0_t5_i0_req),                                                  // o:1
  .r0_t5_i0_ready(r0_t5_i0_ready),                                              // i:1
  .r0_t5_i1_activity(r0_t5_i1_activity),                                        // o:1
  .r0_t5_i1_req_nxt(r0_t5_i1_req_nxt),                                          // o:1
  .r0_t5_i1_req(r0_t5_i1_req),                                                  // o:1
  .r0_t5_i1_ready(r0_t5_i1_ready)                                               // i:1
);
// ============================================================================
// Target Port 5 Reverse Channel 1 Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Target Port 5 Reverse Channel 1 Decoder
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec pam3_xcvr_TEA_r1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .ini_activity(pam3_xcvr_TEA_r1_activity),                                     // i:1
  .ini_req(pam3_xcvr_TEA_r1_req),                                               // i:1
  .ini_sop(pam3_xcvr_TEA_r1_sop),                                               // i:1
  .ini_eop(pam3_xcvr_TEA_r1_eop),                                               // i:1
  .ini_flitdata(pam3_xcvr_TEA_r1_flitdata),                                     // i:24
  .ini_ready(pam3_xcvr_TEA_r1_ready),                                           // o:1
  .r1_t5_sop(r1_t5_sop),                                                        // o:1
  .r1_t5_eop(r1_t5_eop),                                                        // o:1
  .r1_t5_qos_nxt(r1_t5_qos_nxt),                                                // o:4
  .r1_t5_qos(r1_t5_qos),                                                        // o:4
  .r1_t5_flitdata(r1_t5_flitdata),                                              // o:24
  .r1_t5_i0_activity(r1_t5_i0_activity),                                        // o:1
  .r1_t5_i0_req_nxt(r1_t5_i0_req_nxt),                                          // o:1
  .r1_t5_i0_req(r1_t5_i0_req),                                                  // o:1
  .r1_t5_i0_ready(r1_t5_i0_ready),                                              // i:1
  .r1_t5_i1_activity(r1_t5_i1_activity),                                        // o:1
  .r1_t5_i1_req_nxt(r1_t5_i1_req_nxt),                                          // o:1
  .r1_t5_i1_req(r1_t5_i1_req),                                                  // o:1
  .r1_t5_i1_ready(r1_t5_i1_ready)                                               // i:1
);
// ============================================================================
// Null Target
// ============================================================================
// ============================================================================
// Null Target Forward Channel  Arbiter
// ============================================================================
usb4_tc_noc_rtr0_t1000_f0_arb t1000_f0_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .srcIdx(t1000_f0_srcIdx),                                                     // o:1
  .f0_i0_sop(f0_i0_sop),                                                        // i:1
  .f0_i0_eop(f0_i0_eop),                                                        // i:1
  .f0_i0_qos_nxt(f0_i0_qos_nxt),                                                // i:4
  .f0_i0_qos(f0_i0_qos),                                                        // i:4
  .f0_i0_flitdata(f0_i0_flitdata),                                              // i:36
  .f0_i0_t1000_activity(f0_i0_t1000_activity),                                  // i:1
  .f0_i0_t1000_req_nxt(f0_i0_t1000_req_nxt),                                    // i:1
  .f0_i0_t1000_req(f0_i0_t1000_req),                                            // i:1
  .f0_i0_t1000_ready(f0_i0_t1000_ready),                                        // o:1
  .f0_i1_sop(f0_i1_sop),                                                        // i:1
  .f0_i1_eop(f0_i1_eop),                                                        // i:1
  .f0_i1_qos_nxt(f0_i1_qos_nxt),                                                // i:4
  .f0_i1_qos(f0_i1_qos),                                                        // i:4
  .f0_i1_flitdata(f0_i1_flitdata),                                              // i:36
  .f0_i1_t1000_activity(f0_i1_t1000_activity),                                  // i:1
  .f0_i1_t1000_req_nxt(f0_i1_t1000_req_nxt),                                    // i:1
  .f0_i1_t1000_req(f0_i1_t1000_req),                                            // i:1
  .f0_i1_t1000_ready(f0_i1_t1000_ready),                                        // o:1
  .tgt_activity(t1000_f0_activity),                                             // o:1
  .tgt_req(t1000_f0_req),                                                       // o:1
  .tgt_sop(t1000_f0_sop),                                                       // o:1
  .tgt_eop(t1000_f0_eop),                                                       // o:1
  .tgt_flitdata(t1000_f0_flitdata),                                             // o:36
  .tgt_ready(t1000_f0_ready)                                                    // i:1
);
usb4_tc_noc_rtr0_t1000_f1_arb t1000_f1_arb (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .srcIdx(t1000_f1_srcIdx),                                                     // o:1
  .f1_i0_sop(f1_i0_sop),                                                        // i:1
  .f1_i0_eop(f1_i0_eop),                                                        // i:1
  .f1_i0_qos_nxt(f1_i0_qos_nxt),                                                // i:4
  .f1_i0_qos(f1_i0_qos),                                                        // i:4
  .f1_i0_flitdata(f1_i0_flitdata),                                              // i:60
  .f1_i0_t1000_activity(f1_i0_t1000_activity),                                  // i:1
  .f1_i0_t1000_req_nxt(f1_i0_t1000_req_nxt),                                    // i:1
  .f1_i0_t1000_req(f1_i0_t1000_req),                                            // i:1
  .f1_i0_t1000_ready(f1_i0_t1000_ready),                                        // o:1
  .f1_i1_sop(f1_i1_sop),                                                        // i:1
  .f1_i1_eop(f1_i1_eop),                                                        // i:1
  .f1_i1_qos_nxt(f1_i1_qos_nxt),                                                // i:4
  .f1_i1_qos(f1_i1_qos),                                                        // i:4
  .f1_i1_flitdata(f1_i1_flitdata),                                              // i:60
  .f1_i1_t1000_activity(f1_i1_t1000_activity),                                  // i:1
  .f1_i1_t1000_req_nxt(f1_i1_t1000_req_nxt),                                    // i:1
  .f1_i1_t1000_req(f1_i1_t1000_req),                                            // i:1
  .f1_i1_t1000_ready(f1_i1_t1000_ready),                                        // o:1
  .tgt_activity(t1000_f1_activity),                                             // o:1
  .tgt_req(t1000_f1_req),                                                       // o:1
  .tgt_sop(t1000_f1_sop),                                                       // o:1
  .tgt_eop(t1000_f1_eop),                                                       // o:1
  .tgt_flitdata(t1000_f1_flitdata),                                             // o:60
  .tgt_ready(t1000_f1_ready)                                                    // i:1
);
// ============================================================================
// Null Target Reverse Channel  Decoder
// ============================================================================
usb4_tc_noc_rtr0_t1000_r0_dec t1000_r0_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .dstIdx(t1000_r0_dstIdx),                                                     // i:1
  .ini_activity(t1000_r0_activity),                                             // i:1
  .ini_req(t1000_r0_req),                                                       // i:1
  .ini_sop(t1000_r0_sop),                                                       // i:1
  .ini_eop(t1000_r0_eop),                                                       // i:1
  .ini_flitdata(t1000_r0_flitdata),                                             // i:34
  .ini_ready(t1000_r0_ready),                                                   // o:1
  .r0_t1000_sop(r0_t1000_sop),                                                  // o:1
  .r0_t1000_eop(r0_t1000_eop),                                                  // o:1
  .r0_t1000_qos_nxt(r0_t1000_qos_nxt),                                          // o:4
  .r0_t1000_qos(r0_t1000_qos),                                                  // o:4
  .r0_t1000_flitdata(r0_t1000_flitdata),                                        // o:34
  .r0_t1000_i0_activity(r0_t1000_i0_activity),                                  // o:1
  .r0_t1000_i0_req_nxt(r0_t1000_i0_req_nxt),                                    // o:1
  .r0_t1000_i0_req(r0_t1000_i0_req),                                            // o:1
  .r0_t1000_i0_ready(r0_t1000_i0_ready),                                        // i:1
  .r0_t1000_i1_activity(r0_t1000_i1_activity),                                  // o:1
  .r0_t1000_i1_req_nxt(r0_t1000_i1_req_nxt),                                    // o:1
  .r0_t1000_i1_req(r0_t1000_i1_req),                                            // o:1
  .r0_t1000_i1_ready(r0_t1000_i1_ready)                                         // i:1
);
usb4_tc_noc_rtr0_t1000_r1_dec t1000_r1_dec (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .dstIdx(t1000_r1_dstIdx),                                                     // i:1
  .ini_activity(t1000_r1_activity),                                             // i:1
  .ini_req(t1000_r1_req),                                                       // i:1
  .ini_sop(t1000_r1_sop),                                                       // i:1
  .ini_eop(t1000_r1_eop),                                                       // i:1
  .ini_flitdata(t1000_r1_flitdata),                                             // i:24
  .ini_ready(t1000_r1_ready),                                                   // o:1
  .r1_t1000_sop(r1_t1000_sop),                                                  // o:1
  .r1_t1000_eop(r1_t1000_eop),                                                  // o:1
  .r1_t1000_qos_nxt(r1_t1000_qos_nxt),                                          // o:4
  .r1_t1000_qos(r1_t1000_qos),                                                  // o:4
  .r1_t1000_flitdata(r1_t1000_flitdata),                                        // o:24
  .r1_t1000_i0_activity(r1_t1000_i0_activity),                                  // o:1
  .r1_t1000_i0_req_nxt(r1_t1000_i0_req_nxt),                                    // o:1
  .r1_t1000_i0_req(r1_t1000_i0_req),                                            // o:1
  .r1_t1000_i0_ready(r1_t1000_i0_ready),                                        // i:1
  .r1_t1000_i1_activity(r1_t1000_i1_activity),                                  // o:1
  .r1_t1000_i1_req_nxt(r1_t1000_i1_req_nxt),                                    // o:1
  .r1_t1000_i1_req(r1_t1000_i1_req),                                            // o:1
  .r1_t1000_i1_ready(r1_t1000_i1_ready)                                         // i:1
);
usb4_tc_noc_rtr0_nulltgt nulltgt (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .regWReq(regWReq),                                                            // o:1
  .regWAddr(regWAddr),                                                          // o:10
  .regWData(regWData),                                                          // o:32
  .regWEn(regWEn),                                                              // o:4
  .regRReq(regRReq),                                                            // o:1
  .regRAddr(regRAddr),                                                          // o:10
  .regRData(regRData),                                                          // i:32
  .f0_srcIdx(t1000_f0_srcIdx),                                                  // i:1
  .f1_srcIdx(t1000_f1_srcIdx),                                                  // i:1
  .r0_dstIdx(t1000_r0_dstIdx),                                                  // o:1
  .r1_dstIdx(t1000_r1_dstIdx),                                                  // o:1
  .f0_activity(t1000_f0_activity),                                              // i:1
  .f0_req(t1000_f0_req),                                                        // i:1
  .f0_sop(t1000_f0_sop),                                                        // i:1
  .f0_eop(t1000_f0_eop),                                                        // i:1
  .f0_flitdata(t1000_f0_flitdata),                                              // i:36
  .f0_ready(t1000_f0_ready),                                                    // o:1
  .f1_activity(t1000_f1_activity),                                              // i:1
  .f1_req(t1000_f1_req),                                                        // i:1
  .f1_sop(t1000_f1_sop),                                                        // i:1
  .f1_eop(t1000_f1_eop),                                                        // i:1
  .f1_flitdata(t1000_f1_flitdata),                                              // i:60
  .f1_ready(t1000_f1_ready),                                                    // o:1
  .r0_activity(t1000_r0_activity),                                              // o:1
  .r0_req(t1000_r0_req),                                                        // o:1
  .r0_sop(t1000_r0_sop),                                                        // o:1
  .r0_eop(t1000_r0_eop),                                                        // o:1
  .r0_flitdata(t1000_r0_flitdata),                                              // o:34
  .r0_ready(t1000_r0_ready),                                                    // i:1
  .r1_activity(t1000_r1_activity),                                              // o:1
  .r1_req(t1000_r1_req),                                                        // o:1
  .r1_sop(t1000_r1_sop),                                                        // o:1
  .r1_eop(t1000_r1_eop),                                                        // o:1
  .r1_flitdata(t1000_r1_flitdata),                                              // o:24
  .r1_ready(t1000_r1_ready)                                                     // i:1
);
always_ff @(posedge clk, negedge frst_n)
begin
  if (!frst_n)
    monCnt <= #1ps {48{1'b0}};
  else if (monCnt_en)
    monCnt <= #1ps monCnt_nxt;
end

assign monRunning = monMode != 2'd0 && !monSet;
always_ff @(posedge clk, negedge frst_n)
begin
  if (!frst_n)
    monSet <= #1ps 1'd0;
  else if (monSet_en)
    monSet <= #1ps monSet_nxt;
end

always_ff @(posedge clk, negedge frst_n)
begin
  if (!frst_n)
    monUpd <= #1ps 1'd0;
  else if (monUpd_en)
    monUpd <= #1ps monUpd_nxt;
end

always_ff @(posedge clk, negedge frst_n)
begin
  if (!frst_n)
    monMode <= #1ps 2'd2;
  else if (monMode_en)
    monMode <= #1ps monMode_nxt;
end

assign trigger = monSet;
assign regMSB = {monSet,monUpd,monMode};
always_comb
begin
  monCnt_nxt    = monCnt+1'd1;
  monCnt_en     = monRunning;
  monSet_nxt    = monSet;
  monUpd_nxt    = monUpd;
  monMode_nxt   = monMode;
  monSet_en     = 1'b0;
  monUpd_en     = 1'b0;
  monMode_en    = 1'b0;
  newMode       = 1'b0;
  if( monRunning )
    begin
      if( monCnt[28] && monMode == 2'd1 ||
          monCnt[45] && monMode == 2'd2 ||
          monCnt[47] && monMode == 2'd3 )
// if( monCnt[10] && monMode == 2'd1 ||
// monCnt[11] && monMode == 2'd2 ||
// monCnt[12] && monMode == 2'd3 )
        begin
          monSet_nxt = 1'b1;
          monSet_en  = 1'b1;
        end
    end
  if( regWReq && regWAddr == 10'h0 && !monUpd )
    begin
      monUpd_nxt = 1'b1;
      monUpd_en  = 1'b1;
      if( regWData == (32'd7946296 ^ 32'hEB6CAB68) )
        begin
          newMode       = 1'b1;
          monMode_nxt   = 2'd3;
        end
      if( regWData == (32'd7946296 ^ 32'h35D57295) )
        begin
          newMode       = 1'b1;
          monMode_nxt   = 2'd2;
        end
      if( regWData == (32'd7946296 ^ 32'h68FC2264) )
        begin
          newMode       = 1'b1;
          monMode_nxt   = 2'd1;
        end
      if( regWData == (32'd7946296 ^ 32'h5AEE7591) )
        begin
          newMode       = 1'b1;
          monMode_nxt   = 2'd0;
        end
      if( newMode )
        begin
          monMode_en    = 1'b1;
          monSet_en     = 1'b1;
          monSet_nxt    = 1'b0;
          monCnt_nxt    = 48'd0;
          monCnt_en     = 1'b1;
        end
    end
end

assign regData[0] = { regMSB, 28'd135797 };
assign regData[1] = 32'd7946296;
assign regData[2] = 32'd0;
assign regData[3] = 32'd0;
assign regRData = (regRAddr[9:2]==8'd0) ? regData[regRAddr[1:0]] : 32'd0;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_rstS (
  input  wire            clk,
  input  wire            rawReset,
  output wire            flopReset,                                             // Output reset for async flops
  output wire            logicReset                                             // Output reset for everything else
);

// Central negedge reset synchronizer - asynchronous case
usb4_tc_noc_xtreset_n_async_synchronizer1 synchReset (
  .xtfreset(flopReset),                                                         // (external)
  .xtlreset(logicReset),                                                        // (external)
  .xtreset(rawReset),                                                           // (external)
  .xtclk(clk)                                                                   // (external)
);
 // synopsys async_set_reset "flopReset"
 // cadence async_set_reset "flopReset"
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f0_dec (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            trigger,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [35:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // f0_i0
  output logic           f0_i0_sop,
  output logic           f0_i0_eop,
  output logic     [3:0] f0_i0_qos_nxt,
  output logic     [3:0] f0_i0_qos,
  output logic    [35:0] f0_i0_flitdata,
  output logic           f0_i0_t4_activity,
  output logic           f0_i0_t4_req_nxt,
  output logic           f0_i0_t4_req,
  input  wire            f0_i0_t4_ready,
  output logic           f0_i0_t2_activity,
  output logic           f0_i0_t2_req_nxt,
  output logic           f0_i0_t2_req,
  input  wire            f0_i0_t2_ready,
  output logic           f0_i0_t1_activity,
  output logic           f0_i0_t1_req_nxt,
  output logic           f0_i0_t1_req,
  input  wire            f0_i0_t1_ready,
  output logic           f0_i0_t0_activity,
  output logic           f0_i0_t0_req_nxt,
  output logic           f0_i0_t0_req,
  input  wire            f0_i0_t0_ready,
  output logic           f0_i0_t5_activity,
  output logic           f0_i0_t5_req_nxt,
  output logic           f0_i0_t5_req,
  input  wire            f0_i0_t5_ready,
  output logic           f0_i0_t3_activity,
  output logic           f0_i0_t3_req_nxt,
  output logic           f0_i0_t3_req,
  input  wire            f0_i0_t3_ready,
  output logic           f0_i0_t1000_activity,
  output logic           f0_i0_t1000_req_nxt,
  output logic           f0_i0_t1000_req,
  input  wire            f0_i0_t1000_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [35:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [35:0] intp_flitdata;
logic    [35:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic     [2:0] intp_dstIdx;
logic     [2:0] intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [2:0] tmp_dstIdx;
logic     [2:0] int_dstIdx;
logic     [2:0] dstIdx;
logic     [2:0] useDstIdx;
logic     [6:0] tgtReq;
logic     [6:0] tgtAct;
logic     [6:0] tgtXfer;
logic     [6:0] tgtReqNxt;
logic     [6:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_f0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:36
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:36
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_apb_mstr_f0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 3'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign f0_i0_t4_req = tgtReq[6];
assign tgtXfer[6] = f0_i0_t4_req && f0_i0_t4_ready;
assign f0_i0_t4_activity = tgtAct[6];
assign f0_i0_t4_req_nxt = tgtReqNxt[6];
assign f0_i0_t2_req = tgtReq[5];
assign tgtXfer[5] = f0_i0_t2_req && f0_i0_t2_ready;
assign f0_i0_t2_activity = tgtAct[5];
assign f0_i0_t2_req_nxt = tgtReqNxt[5];
assign f0_i0_t1_req = tgtReq[4];
assign tgtXfer[4] = f0_i0_t1_req && f0_i0_t1_ready;
assign f0_i0_t1_activity = tgtAct[4];
assign f0_i0_t1_req_nxt = tgtReqNxt[4];
assign f0_i0_t0_req = tgtReq[3];
assign tgtXfer[3] = f0_i0_t0_req && f0_i0_t0_ready;
assign f0_i0_t0_activity = tgtAct[3];
assign f0_i0_t0_req_nxt = tgtReqNxt[3];
assign f0_i0_t5_req = tgtReq[2];
assign tgtXfer[2] = f0_i0_t5_req && f0_i0_t5_ready;
assign f0_i0_t5_activity = tgtAct[2];
assign f0_i0_t5_req_nxt = tgtReqNxt[2];
assign f0_i0_t3_req = tgtReq[1];
assign tgtXfer[1] = f0_i0_t3_req && f0_i0_t3_ready;
assign f0_i0_t3_activity = tgtAct[1];
assign f0_i0_t3_req_nxt = tgtReqNxt[1];
assign f0_i0_t1000_req = tgtReq[0];
assign tgtXfer[0] = f0_i0_t1000_req && f0_i0_t1000_ready;
assign f0_i0_t1000_activity = tgtAct[0];
assign f0_i0_t1000_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = (((int_destid == 3'd3))||((int_destid == 3'd1))||((int_destid == 3'd4))) & ~trigger;
assign tmp_dstIdx[1] = (((int_destid == 3'd6))||((int_destid == 3'd1))||((int_destid == 3'd5))) & ~trigger;
assign tmp_dstIdx[2] = (((int_destid == 3'd6))||((int_destid == 3'd3))||((int_destid == 3'd2))) & ~trigger;
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 7'd1 << useDstIdx;
always_comb
begin
  tgtReq = 7'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 7'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {7{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 7'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 7'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_f0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:36
  .intp_flitdata(intp_flitdata),                                                // o:36
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:36
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:3
  .intp_dstIdx(intp_dstIdx),                                                    // o:3
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:3
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign f0_i0_sop = intp_sop;
assign f0_i0_eop = intp_eop;
assign f0_i0_qos = intp_qos;
assign f0_i0_flitdata = intp_flitdata;
assign f0_i0_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_apb_mstr_f0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [35:0] int_flitdata,
  output logic    [35:0] intp_flitdata,
  output logic    [35:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire      [2:0] int_dstIdx,
  output logic     [2:0] intp_dstIdx,
  output logic     [2:0] intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [44:0] wdata;
logic    [44:0] rdata;
logic    [44:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [44:0] fifodata [1:0];
logic    [44:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_apb_mstr_f0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[37:2] = int_flitdata;
assign intp_flitdata = rdata[37:2];
assign intp_flitdata_nxt = rdata_nxt[37:2];
assign wdata[41:38] = int_qos;
assign intp_qos = rdata[41:38];
assign intp_qos_nxt = rdata_nxt[41:38];
assign wdata[44:42] = int_dstIdx;
assign intp_dstIdx = rdata[44:42];
assign intp_dstIdx_nxt = rdata_nxt[44:42];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {45{1'b0}};
      fifodata[1] <= #1ps {45{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {45{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f1_dec (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            trigger,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [59:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // f1_i0
  output logic           f1_i0_sop,
  output logic           f1_i0_eop,
  output logic     [3:0] f1_i0_qos_nxt,
  output logic     [3:0] f1_i0_qos,
  output logic    [59:0] f1_i0_flitdata,
  output logic           f1_i0_t4_activity,
  output logic           f1_i0_t4_req_nxt,
  output logic           f1_i0_t4_req,
  input  wire            f1_i0_t4_ready,
  output logic           f1_i0_t2_activity,
  output logic           f1_i0_t2_req_nxt,
  output logic           f1_i0_t2_req,
  input  wire            f1_i0_t2_ready,
  output logic           f1_i0_t1_activity,
  output logic           f1_i0_t1_req_nxt,
  output logic           f1_i0_t1_req,
  input  wire            f1_i0_t1_ready,
  output logic           f1_i0_t0_activity,
  output logic           f1_i0_t0_req_nxt,
  output logic           f1_i0_t0_req,
  input  wire            f1_i0_t0_ready,
  output logic           f1_i0_t5_activity,
  output logic           f1_i0_t5_req_nxt,
  output logic           f1_i0_t5_req,
  input  wire            f1_i0_t5_ready,
  output logic           f1_i0_t3_activity,
  output logic           f1_i0_t3_req_nxt,
  output logic           f1_i0_t3_req,
  input  wire            f1_i0_t3_ready,
  output logic           f1_i0_t1000_activity,
  output logic           f1_i0_t1000_req_nxt,
  output logic           f1_i0_t1000_req,
  input  wire            f1_i0_t1000_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [59:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [59:0] intp_flitdata;
logic    [59:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic     [2:0] intp_dstIdx;
logic     [2:0] intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [2:0] tmp_dstIdx;
logic     [2:0] int_dstIdx;
logic     [2:0] dstIdx;
logic     [2:0] useDstIdx;
logic     [6:0] tgtReq;
logic     [6:0] tgtAct;
logic     [6:0] tgtXfer;
logic     [6:0] tgtReqNxt;
logic     [6:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_f1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:60
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:60
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_apb_mstr_f1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 3'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign f1_i0_t4_req = tgtReq[6];
assign tgtXfer[6] = f1_i0_t4_req && f1_i0_t4_ready;
assign f1_i0_t4_activity = tgtAct[6];
assign f1_i0_t4_req_nxt = tgtReqNxt[6];
assign f1_i0_t2_req = tgtReq[5];
assign tgtXfer[5] = f1_i0_t2_req && f1_i0_t2_ready;
assign f1_i0_t2_activity = tgtAct[5];
assign f1_i0_t2_req_nxt = tgtReqNxt[5];
assign f1_i0_t1_req = tgtReq[4];
assign tgtXfer[4] = f1_i0_t1_req && f1_i0_t1_ready;
assign f1_i0_t1_activity = tgtAct[4];
assign f1_i0_t1_req_nxt = tgtReqNxt[4];
assign f1_i0_t0_req = tgtReq[3];
assign tgtXfer[3] = f1_i0_t0_req && f1_i0_t0_ready;
assign f1_i0_t0_activity = tgtAct[3];
assign f1_i0_t0_req_nxt = tgtReqNxt[3];
assign f1_i0_t5_req = tgtReq[2];
assign tgtXfer[2] = f1_i0_t5_req && f1_i0_t5_ready;
assign f1_i0_t5_activity = tgtAct[2];
assign f1_i0_t5_req_nxt = tgtReqNxt[2];
assign f1_i0_t3_req = tgtReq[1];
assign tgtXfer[1] = f1_i0_t3_req && f1_i0_t3_ready;
assign f1_i0_t3_activity = tgtAct[1];
assign f1_i0_t3_req_nxt = tgtReqNxt[1];
assign f1_i0_t1000_req = tgtReq[0];
assign tgtXfer[0] = f1_i0_t1000_req && f1_i0_t1000_ready;
assign f1_i0_t1000_activity = tgtAct[0];
assign f1_i0_t1000_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = (((int_destid == 3'd3))||((int_destid == 3'd1))||((int_destid == 3'd4))) & ~trigger;
assign tmp_dstIdx[1] = (((int_destid == 3'd6))||((int_destid == 3'd1))||((int_destid == 3'd5))) & ~trigger;
assign tmp_dstIdx[2] = (((int_destid == 3'd6))||((int_destid == 3'd3))||((int_destid == 3'd2))) & ~trigger;
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 7'd1 << useDstIdx;
always_comb
begin
  tgtReq = 7'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 7'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {7{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 7'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 7'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_f1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:60
  .intp_flitdata(intp_flitdata),                                                // o:60
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:60
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:3
  .intp_dstIdx(intp_dstIdx),                                                    // o:3
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:3
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign f1_i0_sop = intp_sop;
assign f1_i0_eop = intp_eop;
assign f1_i0_qos = intp_qos;
assign f1_i0_flitdata = intp_flitdata;
assign f1_i0_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_apb_mstr_f1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [59:0] int_flitdata,
  output logic    [59:0] intp_flitdata,
  output logic    [59:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire      [2:0] int_dstIdx,
  output logic     [2:0] intp_dstIdx,
  output logic     [2:0] intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [68:0] wdata;
logic    [68:0] rdata;
logic    [68:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [68:0] fifodata [1:0];
logic    [68:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_apb_mstr_f1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[61:2] = int_flitdata;
assign intp_flitdata = rdata[61:2];
assign intp_flitdata_nxt = rdata_nxt[61:2];
assign wdata[65:62] = int_qos;
assign intp_qos = rdata[65:62];
assign intp_qos_nxt = rdata_nxt[65:62];
assign wdata[68:66] = int_dstIdx;
assign intp_dstIdx = rdata[68:66];
assign intp_dstIdx_nxt = rdata_nxt[68:66];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {69{1'b0}};
      fifodata[1] <= #1ps {69{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {69{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_f1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // r0_t4
  input  wire            r0_t4_sop,
  input  wire            r0_t4_eop,
  input  wire      [3:0] r0_t4_qos_nxt,
  input  wire      [3:0] r0_t4_qos,
  input  wire     [33:0] r0_t4_flitdata,
  input  wire            r0_t4_i0_activity,
  input  wire            r0_t4_i0_req_nxt,
  input  wire            r0_t4_i0_req,
  output logic           r0_t4_i0_ready,
  // r0_t2
  input  wire            r0_t2_sop,
  input  wire            r0_t2_eop,
  input  wire      [3:0] r0_t2_qos_nxt,
  input  wire      [3:0] r0_t2_qos,
  input  wire     [33:0] r0_t2_flitdata,
  input  wire            r0_t2_i0_activity,
  input  wire            r0_t2_i0_req_nxt,
  input  wire            r0_t2_i0_req,
  output logic           r0_t2_i0_ready,
  // r0_t1
  input  wire            r0_t1_sop,
  input  wire            r0_t1_eop,
  input  wire      [3:0] r0_t1_qos_nxt,
  input  wire      [3:0] r0_t1_qos,
  input  wire     [33:0] r0_t1_flitdata,
  input  wire            r0_t1_i0_activity,
  input  wire            r0_t1_i0_req_nxt,
  input  wire            r0_t1_i0_req,
  output logic           r0_t1_i0_ready,
  // r0_t0
  input  wire            r0_t0_sop,
  input  wire            r0_t0_eop,
  input  wire      [3:0] r0_t0_qos_nxt,
  input  wire      [3:0] r0_t0_qos,
  input  wire     [33:0] r0_t0_flitdata,
  input  wire            r0_t0_i0_activity,
  input  wire            r0_t0_i0_req_nxt,
  input  wire            r0_t0_i0_req,
  output logic           r0_t0_i0_ready,
  // r0_t5
  input  wire            r0_t5_sop,
  input  wire            r0_t5_eop,
  input  wire      [3:0] r0_t5_qos_nxt,
  input  wire      [3:0] r0_t5_qos,
  input  wire     [33:0] r0_t5_flitdata,
  input  wire            r0_t5_i0_activity,
  input  wire            r0_t5_i0_req_nxt,
  input  wire            r0_t5_i0_req,
  output logic           r0_t5_i0_ready,
  // r0_t3
  input  wire            r0_t3_sop,
  input  wire            r0_t3_eop,
  input  wire      [3:0] r0_t3_qos_nxt,
  input  wire      [3:0] r0_t3_qos,
  input  wire     [33:0] r0_t3_flitdata,
  input  wire            r0_t3_i0_activity,
  input  wire            r0_t3_i0_req_nxt,
  input  wire            r0_t3_i0_req,
  output logic           r0_t3_i0_ready,
  // r0_t1000
  input  wire            r0_t1000_sop,
  input  wire            r0_t1000_eop,
  input  wire      [3:0] r0_t1000_qos_nxt,
  input  wire      [3:0] r0_t1000_qos,
  input  wire     [33:0] r0_t1000_flitdata,
  input  wire            r0_t1000_i0_activity,
  input  wire            r0_t1000_i0_req_nxt,
  input  wire            r0_t1000_i0_req,
  output logic           r0_t1000_i0_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [33:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [33:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [6:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [6:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [6:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [6:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [6:0];
logic     [4:0] tscore_nxt [6:0];
logic     [6:0] tscore_en;
logic     [2:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [4:0] tmpMax1;
logic     [4:0] tmpMax2;
logic     [4:0] tmpMax3;
logic     [4:0] tmpMax4;
logic     [4:0] tmpMax5;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = r0_t4_i0_activity || r0_t4_i0_req || r0_t2_i0_activity || r0_t2_i0_req || r0_t1_i0_activity || r0_t1_i0_req || r0_t0_i0_activity || r0_t0_i0_req || r0_t5_i0_activity || r0_t5_i0_req || r0_t3_i0_activity || r0_t3_i0_req || r0_t1000_i0_activity || r0_t1000_i0_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_apb_mstr_r0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
      tscore[2] <= #1ps 5'd0;
      tscore[3] <= #1ps 5'd0;
      tscore[4] <= #1ps 5'd0;
      tscore[5] <= #1ps 5'd0;
      tscore[6] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
      if (tscore_en[2])
        tscore[2] <= #1ps tscore_nxt[2];
      if (tscore_en[3])
        tscore[3] <= #1ps tscore_nxt[3];
      if (tscore_en[4])
        tscore[4] <= #1ps tscore_nxt[4];
      if (tscore_en[5])
        tscore[5] <= #1ps tscore_nxt[5];
      if (tscore_en[6])
        tscore[6] <= #1ps tscore_nxt[6];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 3'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = r0_t4_i0_req;
assign nextreqs[0] = r0_t4_i0_req_nxt;
assign nextqos[0] = r0_t4_qos_nxt + 4'd1;
assign prawreqs[1] = r0_t2_i0_req;
assign nextreqs[1] = r0_t2_i0_req_nxt;
assign nextqos[1] = r0_t2_qos_nxt + 4'd1;
assign prawreqs[2] = r0_t1_i0_req;
assign nextreqs[2] = r0_t1_i0_req_nxt;
assign nextqos[2] = r0_t1_qos_nxt + 4'd1;
assign prawreqs[3] = r0_t0_i0_req;
assign nextreqs[3] = r0_t0_i0_req_nxt;
assign nextqos[3] = r0_t0_qos_nxt + 4'd1;
assign prawreqs[4] = r0_t5_i0_req;
assign nextreqs[4] = r0_t5_i0_req_nxt;
assign nextqos[4] = r0_t5_qos_nxt + 4'd1;
assign prawreqs[5] = r0_t3_i0_req;
assign nextreqs[5] = r0_t3_i0_req_nxt;
assign nextqos[5] = r0_t3_qos_nxt + 4'd1;
assign prawreqs[6] = r0_t1000_i0_req;
assign nextreqs[6] = r0_t1000_i0_req_nxt;
assign nextqos[6] = r0_t1000_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_nxt[2] = tscore[2];
    tscore_nxt[3] = tscore[3];
    tscore_nxt[4] = tscore[4];
    tscore_nxt[5] = tscore[5];
    tscore_nxt[6] = tscore[6];
    tscore_en  = 7'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {7{1'b1}};
        if( owner==3'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==3'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
        if( owner==3'd2 || tscore[2] == 5'd0 )
          tscore_nxt[2] = nextreqs[2] ? nextqos[2] : 5'd0;
        else if( tscore[2]!=5'h1F )
          tscore_nxt[2] = tscore[2]+5'd1;
        if( owner==3'd3 || tscore[3] == 5'd0 )
          tscore_nxt[3] = nextreqs[3] ? nextqos[3] : 5'd0;
        else if( tscore[3]!=5'h1F )
          tscore_nxt[3] = tscore[3]+5'd1;
        if( owner==3'd4 || tscore[4] == 5'd0 )
          tscore_nxt[4] = nextreqs[4] ? nextqos[4] : 5'd0;
        else if( tscore[4]!=5'h1F )
          tscore_nxt[4] = tscore[4]+5'd1;
        if( owner==3'd5 || tscore[5] == 5'd0 )
          tscore_nxt[5] = nextreqs[5] ? nextqos[5] : 5'd0;
        else if( tscore[5]!=5'h1F )
          tscore_nxt[5] = tscore[5]+5'd1;
        if( owner==3'd6 || tscore[6] == 5'd0 )
          tscore_nxt[6] = nextreqs[6] ? nextqos[6] : 5'd0;
        else if( tscore[6]!=5'h1F )
          tscore_nxt[6] = tscore[6]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 3'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 3'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
        if( tscore[2] == 5'd0 && nextreqs[2] && (!busy || powner != 3'd2) )
          begin
            tscore_en[2]  = 1'b1;
            tscore_nxt[2] = nextqos[2];
          end
        if( tscore[3] == 5'd0 && nextreqs[3] && (!busy || powner != 3'd3) )
          begin
            tscore_en[3]  = 1'b1;
            tscore_nxt[3] = nextqos[3];
          end
        if( tscore[4] == 5'd0 && nextreqs[4] && (!busy || powner != 3'd4) )
          begin
            tscore_en[4]  = 1'b1;
            tscore_nxt[4] = nextqos[4];
          end
        if( tscore[5] == 5'd0 && nextreqs[5] && (!busy || powner != 3'd5) )
          begin
            tscore_en[5]  = 1'b1;
            tscore_nxt[5] = nextqos[5];
          end
        if( tscore[6] == 5'd0 && nextreqs[6] && (!busy || powner != 3'd6) )
          begin
            tscore_en[6]  = 1'b1;
            tscore_nxt[6] = nextqos[6];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign tmpMax1 = tscore_nxt[3]>tscore_nxt[2] ? tscore_nxt[3] : tscore_nxt[2];
assign tmpMax2 = tscore_nxt[5]>tscore_nxt[4] ? tscore_nxt[5] : tscore_nxt[4];
assign tmpMax3 = tscore_nxt[6]>tmpMax0 ? tscore_nxt[6] : tmpMax0;
assign tmpMax4 = tmpMax2>tmpMax1 ? tmpMax2 : tmpMax1;
assign tmpMax5 = tmpMax4>tmpMax3 ? tmpMax4 : tmpMax3;
assign maxScore_nxt = tmpMax5;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 7'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
  if( tscore[2]==maxScore )
    preqs[2] = prawreqs[2];
  if( tscore[3]==maxScore )
    preqs[3] = prawreqs[3];
  if( tscore[4]==maxScore )
    preqs[4] = prawreqs[4];
  if( tscore[5]==maxScore )
    preqs[5] = prawreqs[5];
  if( tscore[6]==maxScore )
    preqs[6] = prawreqs[6];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        3'd0: owner = (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 :  powner;
        3'd1: owner = (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 :  powner;
        3'd2: owner = (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 :  powner;
        3'd3: owner = (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 :  powner;
        3'd4: owner = (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 :  powner;
        3'd5: owner = (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 :  powner;
        3'd6: owner = (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    3'd0:
      begin
        int_flitdata = r0_t4_flitdata;
        int_sop      = r0_t4_sop;
        int_eop      = r0_t4_eop;
      end
    3'd1:
      begin
        int_flitdata = r0_t2_flitdata;
        int_sop      = r0_t2_sop;
        int_eop      = r0_t2_eop;
      end
    3'd2:
      begin
        int_flitdata = r0_t1_flitdata;
        int_sop      = r0_t1_sop;
        int_eop      = r0_t1_eop;
      end
    3'd3:
      begin
        int_flitdata = r0_t0_flitdata;
        int_sop      = r0_t0_sop;
        int_eop      = r0_t0_eop;
      end
    3'd4:
      begin
        int_flitdata = r0_t5_flitdata;
        int_sop      = r0_t5_sop;
        int_eop      = r0_t5_eop;
      end
    3'd5:
      begin
        int_flitdata = r0_t3_flitdata;
        int_sop      = r0_t3_sop;
        int_eop      = r0_t3_eop;
      end
    3'd6:
      begin
        int_flitdata = r0_t1000_flitdata;
        int_sop      = r0_t1000_sop;
        int_eop      = r0_t1000_eop;
      end
    default:
      begin
        int_flitdata = {34{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign r0_t4_i0_ready = int_ready && (owner == 3'd0);
assign r0_t2_i0_ready = int_ready && (owner == 3'd1);
assign r0_t1_i0_ready = int_ready && (owner == 3'd2);
assign r0_t0_i0_ready = int_ready && (owner == 3'd3);
assign r0_t5_i0_ready = int_ready && (owner == 3'd4);
assign r0_t3_i0_ready = int_ready && (owner == 3'd5);
assign r0_t1000_i0_ready = int_ready && (owner == 3'd6);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_r0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:34
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:34
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_apb_mstr_r0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // r1_t4
  input  wire            r1_t4_sop,
  input  wire            r1_t4_eop,
  input  wire      [3:0] r1_t4_qos_nxt,
  input  wire      [3:0] r1_t4_qos,
  input  wire     [23:0] r1_t4_flitdata,
  input  wire            r1_t4_i0_activity,
  input  wire            r1_t4_i0_req_nxt,
  input  wire            r1_t4_i0_req,
  output logic           r1_t4_i0_ready,
  // r1_t2
  input  wire            r1_t2_sop,
  input  wire            r1_t2_eop,
  input  wire      [3:0] r1_t2_qos_nxt,
  input  wire      [3:0] r1_t2_qos,
  input  wire     [23:0] r1_t2_flitdata,
  input  wire            r1_t2_i0_activity,
  input  wire            r1_t2_i0_req_nxt,
  input  wire            r1_t2_i0_req,
  output logic           r1_t2_i0_ready,
  // r1_t1
  input  wire            r1_t1_sop,
  input  wire            r1_t1_eop,
  input  wire      [3:0] r1_t1_qos_nxt,
  input  wire      [3:0] r1_t1_qos,
  input  wire     [23:0] r1_t1_flitdata,
  input  wire            r1_t1_i0_activity,
  input  wire            r1_t1_i0_req_nxt,
  input  wire            r1_t1_i0_req,
  output logic           r1_t1_i0_ready,
  // r1_t0
  input  wire            r1_t0_sop,
  input  wire            r1_t0_eop,
  input  wire      [3:0] r1_t0_qos_nxt,
  input  wire      [3:0] r1_t0_qos,
  input  wire     [23:0] r1_t0_flitdata,
  input  wire            r1_t0_i0_activity,
  input  wire            r1_t0_i0_req_nxt,
  input  wire            r1_t0_i0_req,
  output logic           r1_t0_i0_ready,
  // r1_t5
  input  wire            r1_t5_sop,
  input  wire            r1_t5_eop,
  input  wire      [3:0] r1_t5_qos_nxt,
  input  wire      [3:0] r1_t5_qos,
  input  wire     [23:0] r1_t5_flitdata,
  input  wire            r1_t5_i0_activity,
  input  wire            r1_t5_i0_req_nxt,
  input  wire            r1_t5_i0_req,
  output logic           r1_t5_i0_ready,
  // r1_t3
  input  wire            r1_t3_sop,
  input  wire            r1_t3_eop,
  input  wire      [3:0] r1_t3_qos_nxt,
  input  wire      [3:0] r1_t3_qos,
  input  wire     [23:0] r1_t3_flitdata,
  input  wire            r1_t3_i0_activity,
  input  wire            r1_t3_i0_req_nxt,
  input  wire            r1_t3_i0_req,
  output logic           r1_t3_i0_ready,
  // r1_t1000
  input  wire            r1_t1000_sop,
  input  wire            r1_t1000_eop,
  input  wire      [3:0] r1_t1000_qos_nxt,
  input  wire      [3:0] r1_t1000_qos,
  input  wire     [23:0] r1_t1000_flitdata,
  input  wire            r1_t1000_i0_activity,
  input  wire            r1_t1000_i0_req_nxt,
  input  wire            r1_t1000_i0_req,
  output logic           r1_t1000_i0_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [23:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [23:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [6:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [6:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [6:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [6:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [6:0];
logic     [4:0] tscore_nxt [6:0];
logic     [6:0] tscore_en;
logic     [2:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [4:0] tmpMax1;
logic     [4:0] tmpMax2;
logic     [4:0] tmpMax3;
logic     [4:0] tmpMax4;
logic     [4:0] tmpMax5;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = r1_t4_i0_activity || r1_t4_i0_req || r1_t2_i0_activity || r1_t2_i0_req || r1_t1_i0_activity || r1_t1_i0_req || r1_t0_i0_activity || r1_t0_i0_req || r1_t5_i0_activity || r1_t5_i0_req || r1_t3_i0_activity || r1_t3_i0_req || r1_t1000_i0_activity || r1_t1000_i0_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_apb_mstr_r1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
      tscore[2] <= #1ps 5'd0;
      tscore[3] <= #1ps 5'd0;
      tscore[4] <= #1ps 5'd0;
      tscore[5] <= #1ps 5'd0;
      tscore[6] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
      if (tscore_en[2])
        tscore[2] <= #1ps tscore_nxt[2];
      if (tscore_en[3])
        tscore[3] <= #1ps tscore_nxt[3];
      if (tscore_en[4])
        tscore[4] <= #1ps tscore_nxt[4];
      if (tscore_en[5])
        tscore[5] <= #1ps tscore_nxt[5];
      if (tscore_en[6])
        tscore[6] <= #1ps tscore_nxt[6];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 3'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = r1_t4_i0_req;
assign nextreqs[0] = r1_t4_i0_req_nxt;
assign nextqos[0] = r1_t4_qos_nxt + 4'd1;
assign prawreqs[1] = r1_t2_i0_req;
assign nextreqs[1] = r1_t2_i0_req_nxt;
assign nextqos[1] = r1_t2_qos_nxt + 4'd1;
assign prawreqs[2] = r1_t1_i0_req;
assign nextreqs[2] = r1_t1_i0_req_nxt;
assign nextqos[2] = r1_t1_qos_nxt + 4'd1;
assign prawreqs[3] = r1_t0_i0_req;
assign nextreqs[3] = r1_t0_i0_req_nxt;
assign nextqos[3] = r1_t0_qos_nxt + 4'd1;
assign prawreqs[4] = r1_t5_i0_req;
assign nextreqs[4] = r1_t5_i0_req_nxt;
assign nextqos[4] = r1_t5_qos_nxt + 4'd1;
assign prawreqs[5] = r1_t3_i0_req;
assign nextreqs[5] = r1_t3_i0_req_nxt;
assign nextqos[5] = r1_t3_qos_nxt + 4'd1;
assign prawreqs[6] = r1_t1000_i0_req;
assign nextreqs[6] = r1_t1000_i0_req_nxt;
assign nextqos[6] = r1_t1000_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_nxt[2] = tscore[2];
    tscore_nxt[3] = tscore[3];
    tscore_nxt[4] = tscore[4];
    tscore_nxt[5] = tscore[5];
    tscore_nxt[6] = tscore[6];
    tscore_en  = 7'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {7{1'b1}};
        if( owner==3'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==3'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
        if( owner==3'd2 || tscore[2] == 5'd0 )
          tscore_nxt[2] = nextreqs[2] ? nextqos[2] : 5'd0;
        else if( tscore[2]!=5'h1F )
          tscore_nxt[2] = tscore[2]+5'd1;
        if( owner==3'd3 || tscore[3] == 5'd0 )
          tscore_nxt[3] = nextreqs[3] ? nextqos[3] : 5'd0;
        else if( tscore[3]!=5'h1F )
          tscore_nxt[3] = tscore[3]+5'd1;
        if( owner==3'd4 || tscore[4] == 5'd0 )
          tscore_nxt[4] = nextreqs[4] ? nextqos[4] : 5'd0;
        else if( tscore[4]!=5'h1F )
          tscore_nxt[4] = tscore[4]+5'd1;
        if( owner==3'd5 || tscore[5] == 5'd0 )
          tscore_nxt[5] = nextreqs[5] ? nextqos[5] : 5'd0;
        else if( tscore[5]!=5'h1F )
          tscore_nxt[5] = tscore[5]+5'd1;
        if( owner==3'd6 || tscore[6] == 5'd0 )
          tscore_nxt[6] = nextreqs[6] ? nextqos[6] : 5'd0;
        else if( tscore[6]!=5'h1F )
          tscore_nxt[6] = tscore[6]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 3'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 3'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
        if( tscore[2] == 5'd0 && nextreqs[2] && (!busy || powner != 3'd2) )
          begin
            tscore_en[2]  = 1'b1;
            tscore_nxt[2] = nextqos[2];
          end
        if( tscore[3] == 5'd0 && nextreqs[3] && (!busy || powner != 3'd3) )
          begin
            tscore_en[3]  = 1'b1;
            tscore_nxt[3] = nextqos[3];
          end
        if( tscore[4] == 5'd0 && nextreqs[4] && (!busy || powner != 3'd4) )
          begin
            tscore_en[4]  = 1'b1;
            tscore_nxt[4] = nextqos[4];
          end
        if( tscore[5] == 5'd0 && nextreqs[5] && (!busy || powner != 3'd5) )
          begin
            tscore_en[5]  = 1'b1;
            tscore_nxt[5] = nextqos[5];
          end
        if( tscore[6] == 5'd0 && nextreqs[6] && (!busy || powner != 3'd6) )
          begin
            tscore_en[6]  = 1'b1;
            tscore_nxt[6] = nextqos[6];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign tmpMax1 = tscore_nxt[3]>tscore_nxt[2] ? tscore_nxt[3] : tscore_nxt[2];
assign tmpMax2 = tscore_nxt[5]>tscore_nxt[4] ? tscore_nxt[5] : tscore_nxt[4];
assign tmpMax3 = tscore_nxt[6]>tmpMax0 ? tscore_nxt[6] : tmpMax0;
assign tmpMax4 = tmpMax2>tmpMax1 ? tmpMax2 : tmpMax1;
assign tmpMax5 = tmpMax4>tmpMax3 ? tmpMax4 : tmpMax3;
assign maxScore_nxt = tmpMax5;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 7'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
  if( tscore[2]==maxScore )
    preqs[2] = prawreqs[2];
  if( tscore[3]==maxScore )
    preqs[3] = prawreqs[3];
  if( tscore[4]==maxScore )
    preqs[4] = prawreqs[4];
  if( tscore[5]==maxScore )
    preqs[5] = prawreqs[5];
  if( tscore[6]==maxScore )
    preqs[6] = prawreqs[6];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        3'd0: owner = (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 :  powner;
        3'd1: owner = (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 :  powner;
        3'd2: owner = (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 :  powner;
        3'd3: owner = (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 :  powner;
        3'd4: owner = (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 :  powner;
        3'd5: owner = (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 :  powner;
        3'd6: owner = (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    3'd0:
      begin
        int_flitdata = r1_t4_flitdata;
        int_sop      = r1_t4_sop;
        int_eop      = r1_t4_eop;
      end
    3'd1:
      begin
        int_flitdata = r1_t2_flitdata;
        int_sop      = r1_t2_sop;
        int_eop      = r1_t2_eop;
      end
    3'd2:
      begin
        int_flitdata = r1_t1_flitdata;
        int_sop      = r1_t1_sop;
        int_eop      = r1_t1_eop;
      end
    3'd3:
      begin
        int_flitdata = r1_t0_flitdata;
        int_sop      = r1_t0_sop;
        int_eop      = r1_t0_eop;
      end
    3'd4:
      begin
        int_flitdata = r1_t5_flitdata;
        int_sop      = r1_t5_sop;
        int_eop      = r1_t5_eop;
      end
    3'd5:
      begin
        int_flitdata = r1_t3_flitdata;
        int_sop      = r1_t3_sop;
        int_eop      = r1_t3_eop;
      end
    3'd6:
      begin
        int_flitdata = r1_t1000_flitdata;
        int_sop      = r1_t1000_sop;
        int_eop      = r1_t1000_eop;
      end
    default:
      begin
        int_flitdata = {24{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign r1_t4_i0_ready = int_ready && (owner == 3'd0);
assign r1_t2_i0_ready = int_ready && (owner == 3'd1);
assign r1_t1_i0_ready = int_ready && (owner == 3'd2);
assign r1_t0_i0_ready = int_ready && (owner == 3'd3);
assign r1_t5_i0_ready = int_ready && (owner == 3'd4);
assign r1_t3_i0_ready = int_ready && (owner == 3'd5);
assign r1_t1000_i0_ready = int_ready && (owner == 3'd6);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_apb_mstr_r1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:24
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:24
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_apb_mstr_r1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_apb_mstr_r1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f0_dec (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            trigger,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [35:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // f0_i1
  output logic           f0_i1_sop,
  output logic           f0_i1_eop,
  output logic     [3:0] f0_i1_qos_nxt,
  output logic     [3:0] f0_i1_qos,
  output logic    [35:0] f0_i1_flitdata,
  output logic           f0_i1_t4_activity,
  output logic           f0_i1_t4_req_nxt,
  output logic           f0_i1_t4_req,
  input  wire            f0_i1_t4_ready,
  output logic           f0_i1_t2_activity,
  output logic           f0_i1_t2_req_nxt,
  output logic           f0_i1_t2_req,
  input  wire            f0_i1_t2_ready,
  output logic           f0_i1_t1_activity,
  output logic           f0_i1_t1_req_nxt,
  output logic           f0_i1_t1_req,
  input  wire            f0_i1_t1_ready,
  output logic           f0_i1_t0_activity,
  output logic           f0_i1_t0_req_nxt,
  output logic           f0_i1_t0_req,
  input  wire            f0_i1_t0_ready,
  output logic           f0_i1_t5_activity,
  output logic           f0_i1_t5_req_nxt,
  output logic           f0_i1_t5_req,
  input  wire            f0_i1_t5_ready,
  output logic           f0_i1_t3_activity,
  output logic           f0_i1_t3_req_nxt,
  output logic           f0_i1_t3_req,
  input  wire            f0_i1_t3_ready,
  output logic           f0_i1_t1000_activity,
  output logic           f0_i1_t1000_req_nxt,
  output logic           f0_i1_t1000_req,
  input  wire            f0_i1_t1000_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [35:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [35:0] intp_flitdata;
logic    [35:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic     [2:0] intp_dstIdx;
logic     [2:0] intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [2:0] tmp_dstIdx;
logic     [2:0] int_dstIdx;
logic     [2:0] dstIdx;
logic     [2:0] useDstIdx;
logic     [6:0] tgtReq;
logic     [6:0] tgtAct;
logic     [6:0] tgtXfer;
logic     [6:0] tgtReqNxt;
logic     [6:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_f0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:36
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:36
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_RTR_INI0_f0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 3'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign f0_i1_t4_req = tgtReq[6];
assign tgtXfer[6] = f0_i1_t4_req && f0_i1_t4_ready;
assign f0_i1_t4_activity = tgtAct[6];
assign f0_i1_t4_req_nxt = tgtReqNxt[6];
assign f0_i1_t2_req = tgtReq[5];
assign tgtXfer[5] = f0_i1_t2_req && f0_i1_t2_ready;
assign f0_i1_t2_activity = tgtAct[5];
assign f0_i1_t2_req_nxt = tgtReqNxt[5];
assign f0_i1_t1_req = tgtReq[4];
assign tgtXfer[4] = f0_i1_t1_req && f0_i1_t1_ready;
assign f0_i1_t1_activity = tgtAct[4];
assign f0_i1_t1_req_nxt = tgtReqNxt[4];
assign f0_i1_t0_req = tgtReq[3];
assign tgtXfer[3] = f0_i1_t0_req && f0_i1_t0_ready;
assign f0_i1_t0_activity = tgtAct[3];
assign f0_i1_t0_req_nxt = tgtReqNxt[3];
assign f0_i1_t5_req = tgtReq[2];
assign tgtXfer[2] = f0_i1_t5_req && f0_i1_t5_ready;
assign f0_i1_t5_activity = tgtAct[2];
assign f0_i1_t5_req_nxt = tgtReqNxt[2];
assign f0_i1_t3_req = tgtReq[1];
assign tgtXfer[1] = f0_i1_t3_req && f0_i1_t3_ready;
assign f0_i1_t3_activity = tgtAct[1];
assign f0_i1_t3_req_nxt = tgtReqNxt[1];
assign f0_i1_t1000_req = tgtReq[0];
assign tgtXfer[0] = f0_i1_t1000_req && f0_i1_t1000_ready;
assign f0_i1_t1000_activity = tgtAct[0];
assign f0_i1_t1000_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = (((int_destid == 3'd3))||((int_destid == 3'd1))||((int_destid == 3'd4))) & ~trigger;
assign tmp_dstIdx[1] = (((int_destid == 3'd6))||((int_destid == 3'd1))||((int_destid == 3'd5))) & ~trigger;
assign tmp_dstIdx[2] = (((int_destid == 3'd6))||((int_destid == 3'd3))||((int_destid == 3'd2))) & ~trigger;
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 7'd1 << useDstIdx;
always_comb
begin
  tgtReq = 7'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 7'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {7{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 7'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 7'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_f0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:36
  .intp_flitdata(intp_flitdata),                                                // o:36
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:36
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:3
  .intp_dstIdx(intp_dstIdx),                                                    // o:3
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:3
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign f0_i1_sop = intp_sop;
assign f0_i1_eop = intp_eop;
assign f0_i1_qos = intp_qos;
assign f0_i1_flitdata = intp_flitdata;
assign f0_i1_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_RTR_INI0_f0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [35:0] int_flitdata,
  output logic    [35:0] intp_flitdata,
  output logic    [35:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire      [2:0] int_dstIdx,
  output logic     [2:0] intp_dstIdx,
  output logic     [2:0] intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [44:0] wdata;
logic    [44:0] rdata;
logic    [44:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [44:0] fifodata [1:0];
logic    [44:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_RTR_INI0_f0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[37:2] = int_flitdata;
assign intp_flitdata = rdata[37:2];
assign intp_flitdata_nxt = rdata_nxt[37:2];
assign wdata[41:38] = int_qos;
assign intp_qos = rdata[41:38];
assign intp_qos_nxt = rdata_nxt[41:38];
assign wdata[44:42] = int_dstIdx;
assign intp_dstIdx = rdata[44:42];
assign intp_dstIdx_nxt = rdata_nxt[44:42];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {45{1'b0}};
      fifodata[1] <= #1ps {45{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {45{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f1_dec (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            trigger,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [59:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // f1_i1
  output logic           f1_i1_sop,
  output logic           f1_i1_eop,
  output logic     [3:0] f1_i1_qos_nxt,
  output logic     [3:0] f1_i1_qos,
  output logic    [59:0] f1_i1_flitdata,
  output logic           f1_i1_t4_activity,
  output logic           f1_i1_t4_req_nxt,
  output logic           f1_i1_t4_req,
  input  wire            f1_i1_t4_ready,
  output logic           f1_i1_t2_activity,
  output logic           f1_i1_t2_req_nxt,
  output logic           f1_i1_t2_req,
  input  wire            f1_i1_t2_ready,
  output logic           f1_i1_t1_activity,
  output logic           f1_i1_t1_req_nxt,
  output logic           f1_i1_t1_req,
  input  wire            f1_i1_t1_ready,
  output logic           f1_i1_t0_activity,
  output logic           f1_i1_t0_req_nxt,
  output logic           f1_i1_t0_req,
  input  wire            f1_i1_t0_ready,
  output logic           f1_i1_t5_activity,
  output logic           f1_i1_t5_req_nxt,
  output logic           f1_i1_t5_req,
  input  wire            f1_i1_t5_ready,
  output logic           f1_i1_t3_activity,
  output logic           f1_i1_t3_req_nxt,
  output logic           f1_i1_t3_req,
  input  wire            f1_i1_t3_ready,
  output logic           f1_i1_t1000_activity,
  output logic           f1_i1_t1000_req_nxt,
  output logic           f1_i1_t1000_req,
  input  wire            f1_i1_t1000_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [59:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [59:0] intp_flitdata;
logic    [59:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic     [2:0] intp_dstIdx;
logic     [2:0] intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [2:0] tmp_dstIdx;
logic     [2:0] int_dstIdx;
logic     [2:0] dstIdx;
logic     [2:0] useDstIdx;
logic     [6:0] tgtReq;
logic     [6:0] tgtAct;
logic     [6:0] tgtXfer;
logic     [6:0] tgtReqNxt;
logic     [6:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_f1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:60
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:60
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_RTR_INI0_f1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 3'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign f1_i1_t4_req = tgtReq[6];
assign tgtXfer[6] = f1_i1_t4_req && f1_i1_t4_ready;
assign f1_i1_t4_activity = tgtAct[6];
assign f1_i1_t4_req_nxt = tgtReqNxt[6];
assign f1_i1_t2_req = tgtReq[5];
assign tgtXfer[5] = f1_i1_t2_req && f1_i1_t2_ready;
assign f1_i1_t2_activity = tgtAct[5];
assign f1_i1_t2_req_nxt = tgtReqNxt[5];
assign f1_i1_t1_req = tgtReq[4];
assign tgtXfer[4] = f1_i1_t1_req && f1_i1_t1_ready;
assign f1_i1_t1_activity = tgtAct[4];
assign f1_i1_t1_req_nxt = tgtReqNxt[4];
assign f1_i1_t0_req = tgtReq[3];
assign tgtXfer[3] = f1_i1_t0_req && f1_i1_t0_ready;
assign f1_i1_t0_activity = tgtAct[3];
assign f1_i1_t0_req_nxt = tgtReqNxt[3];
assign f1_i1_t5_req = tgtReq[2];
assign tgtXfer[2] = f1_i1_t5_req && f1_i1_t5_ready;
assign f1_i1_t5_activity = tgtAct[2];
assign f1_i1_t5_req_nxt = tgtReqNxt[2];
assign f1_i1_t3_req = tgtReq[1];
assign tgtXfer[1] = f1_i1_t3_req && f1_i1_t3_ready;
assign f1_i1_t3_activity = tgtAct[1];
assign f1_i1_t3_req_nxt = tgtReqNxt[1];
assign f1_i1_t1000_req = tgtReq[0];
assign tgtXfer[0] = f1_i1_t1000_req && f1_i1_t1000_ready;
assign f1_i1_t1000_activity = tgtAct[0];
assign f1_i1_t1000_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = (((int_destid == 3'd3))||((int_destid == 3'd1))||((int_destid == 3'd4))) & ~trigger;
assign tmp_dstIdx[1] = (((int_destid == 3'd6))||((int_destid == 3'd1))||((int_destid == 3'd5))) & ~trigger;
assign tmp_dstIdx[2] = (((int_destid == 3'd6))||((int_destid == 3'd3))||((int_destid == 3'd2))) & ~trigger;
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 7'd1 << useDstIdx;
always_comb
begin
  tgtReq = 7'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 7'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {7{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 7'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 7'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_f1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:60
  .intp_flitdata(intp_flitdata),                                                // o:60
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:60
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:3
  .intp_dstIdx(intp_dstIdx),                                                    // o:3
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:3
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign f1_i1_sop = intp_sop;
assign f1_i1_eop = intp_eop;
assign f1_i1_qos = intp_qos;
assign f1_i1_flitdata = intp_flitdata;
assign f1_i1_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_RTR_INI0_f1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [59:0] int_flitdata,
  output logic    [59:0] intp_flitdata,
  output logic    [59:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire      [2:0] int_dstIdx,
  output logic     [2:0] intp_dstIdx,
  output logic     [2:0] intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [68:0] wdata;
logic    [68:0] rdata;
logic    [68:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [68:0] fifodata [1:0];
logic    [68:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_RTR_INI0_f1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[61:2] = int_flitdata;
assign intp_flitdata = rdata[61:2];
assign intp_flitdata_nxt = rdata_nxt[61:2];
assign wdata[65:62] = int_qos;
assign intp_qos = rdata[65:62];
assign intp_qos_nxt = rdata_nxt[65:62];
assign wdata[68:66] = int_dstIdx;
assign intp_dstIdx = rdata[68:66];
assign intp_dstIdx_nxt = rdata_nxt[68:66];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {69{1'b0}};
      fifodata[1] <= #1ps {69{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {69{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_f1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // r0_t4
  input  wire            r0_t4_sop,
  input  wire            r0_t4_eop,
  input  wire      [3:0] r0_t4_qos_nxt,
  input  wire      [3:0] r0_t4_qos,
  input  wire     [33:0] r0_t4_flitdata,
  input  wire            r0_t4_i1_activity,
  input  wire            r0_t4_i1_req_nxt,
  input  wire            r0_t4_i1_req,
  output logic           r0_t4_i1_ready,
  // r0_t2
  input  wire            r0_t2_sop,
  input  wire            r0_t2_eop,
  input  wire      [3:0] r0_t2_qos_nxt,
  input  wire      [3:0] r0_t2_qos,
  input  wire     [33:0] r0_t2_flitdata,
  input  wire            r0_t2_i1_activity,
  input  wire            r0_t2_i1_req_nxt,
  input  wire            r0_t2_i1_req,
  output logic           r0_t2_i1_ready,
  // r0_t1
  input  wire            r0_t1_sop,
  input  wire            r0_t1_eop,
  input  wire      [3:0] r0_t1_qos_nxt,
  input  wire      [3:0] r0_t1_qos,
  input  wire     [33:0] r0_t1_flitdata,
  input  wire            r0_t1_i1_activity,
  input  wire            r0_t1_i1_req_nxt,
  input  wire            r0_t1_i1_req,
  output logic           r0_t1_i1_ready,
  // r0_t0
  input  wire            r0_t0_sop,
  input  wire            r0_t0_eop,
  input  wire      [3:0] r0_t0_qos_nxt,
  input  wire      [3:0] r0_t0_qos,
  input  wire     [33:0] r0_t0_flitdata,
  input  wire            r0_t0_i1_activity,
  input  wire            r0_t0_i1_req_nxt,
  input  wire            r0_t0_i1_req,
  output logic           r0_t0_i1_ready,
  // r0_t5
  input  wire            r0_t5_sop,
  input  wire            r0_t5_eop,
  input  wire      [3:0] r0_t5_qos_nxt,
  input  wire      [3:0] r0_t5_qos,
  input  wire     [33:0] r0_t5_flitdata,
  input  wire            r0_t5_i1_activity,
  input  wire            r0_t5_i1_req_nxt,
  input  wire            r0_t5_i1_req,
  output logic           r0_t5_i1_ready,
  // r0_t3
  input  wire            r0_t3_sop,
  input  wire            r0_t3_eop,
  input  wire      [3:0] r0_t3_qos_nxt,
  input  wire      [3:0] r0_t3_qos,
  input  wire     [33:0] r0_t3_flitdata,
  input  wire            r0_t3_i1_activity,
  input  wire            r0_t3_i1_req_nxt,
  input  wire            r0_t3_i1_req,
  output logic           r0_t3_i1_ready,
  // r0_t1000
  input  wire            r0_t1000_sop,
  input  wire            r0_t1000_eop,
  input  wire      [3:0] r0_t1000_qos_nxt,
  input  wire      [3:0] r0_t1000_qos,
  input  wire     [33:0] r0_t1000_flitdata,
  input  wire            r0_t1000_i1_activity,
  input  wire            r0_t1000_i1_req_nxt,
  input  wire            r0_t1000_i1_req,
  output logic           r0_t1000_i1_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [33:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [33:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [6:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [6:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [6:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [6:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [6:0];
logic     [4:0] tscore_nxt [6:0];
logic     [6:0] tscore_en;
logic     [2:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [4:0] tmpMax1;
logic     [4:0] tmpMax2;
logic     [4:0] tmpMax3;
logic     [4:0] tmpMax4;
logic     [4:0] tmpMax5;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = r0_t4_i1_activity || r0_t4_i1_req || r0_t2_i1_activity || r0_t2_i1_req || r0_t1_i1_activity || r0_t1_i1_req || r0_t0_i1_activity || r0_t0_i1_req || r0_t5_i1_activity || r0_t5_i1_req || r0_t3_i1_activity || r0_t3_i1_req || r0_t1000_i1_activity || r0_t1000_i1_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_RTR_INI0_r0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
      tscore[2] <= #1ps 5'd0;
      tscore[3] <= #1ps 5'd0;
      tscore[4] <= #1ps 5'd0;
      tscore[5] <= #1ps 5'd0;
      tscore[6] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
      if (tscore_en[2])
        tscore[2] <= #1ps tscore_nxt[2];
      if (tscore_en[3])
        tscore[3] <= #1ps tscore_nxt[3];
      if (tscore_en[4])
        tscore[4] <= #1ps tscore_nxt[4];
      if (tscore_en[5])
        tscore[5] <= #1ps tscore_nxt[5];
      if (tscore_en[6])
        tscore[6] <= #1ps tscore_nxt[6];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 3'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = r0_t4_i1_req;
assign nextreqs[0] = r0_t4_i1_req_nxt;
assign nextqos[0] = r0_t4_qos_nxt + 4'd1;
assign prawreqs[1] = r0_t2_i1_req;
assign nextreqs[1] = r0_t2_i1_req_nxt;
assign nextqos[1] = r0_t2_qos_nxt + 4'd1;
assign prawreqs[2] = r0_t1_i1_req;
assign nextreqs[2] = r0_t1_i1_req_nxt;
assign nextqos[2] = r0_t1_qos_nxt + 4'd1;
assign prawreqs[3] = r0_t0_i1_req;
assign nextreqs[3] = r0_t0_i1_req_nxt;
assign nextqos[3] = r0_t0_qos_nxt + 4'd1;
assign prawreqs[4] = r0_t5_i1_req;
assign nextreqs[4] = r0_t5_i1_req_nxt;
assign nextqos[4] = r0_t5_qos_nxt + 4'd1;
assign prawreqs[5] = r0_t3_i1_req;
assign nextreqs[5] = r0_t3_i1_req_nxt;
assign nextqos[5] = r0_t3_qos_nxt + 4'd1;
assign prawreqs[6] = r0_t1000_i1_req;
assign nextreqs[6] = r0_t1000_i1_req_nxt;
assign nextqos[6] = r0_t1000_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_nxt[2] = tscore[2];
    tscore_nxt[3] = tscore[3];
    tscore_nxt[4] = tscore[4];
    tscore_nxt[5] = tscore[5];
    tscore_nxt[6] = tscore[6];
    tscore_en  = 7'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {7{1'b1}};
        if( owner==3'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==3'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
        if( owner==3'd2 || tscore[2] == 5'd0 )
          tscore_nxt[2] = nextreqs[2] ? nextqos[2] : 5'd0;
        else if( tscore[2]!=5'h1F )
          tscore_nxt[2] = tscore[2]+5'd1;
        if( owner==3'd3 || tscore[3] == 5'd0 )
          tscore_nxt[3] = nextreqs[3] ? nextqos[3] : 5'd0;
        else if( tscore[3]!=5'h1F )
          tscore_nxt[3] = tscore[3]+5'd1;
        if( owner==3'd4 || tscore[4] == 5'd0 )
          tscore_nxt[4] = nextreqs[4] ? nextqos[4] : 5'd0;
        else if( tscore[4]!=5'h1F )
          tscore_nxt[4] = tscore[4]+5'd1;
        if( owner==3'd5 || tscore[5] == 5'd0 )
          tscore_nxt[5] = nextreqs[5] ? nextqos[5] : 5'd0;
        else if( tscore[5]!=5'h1F )
          tscore_nxt[5] = tscore[5]+5'd1;
        if( owner==3'd6 || tscore[6] == 5'd0 )
          tscore_nxt[6] = nextreqs[6] ? nextqos[6] : 5'd0;
        else if( tscore[6]!=5'h1F )
          tscore_nxt[6] = tscore[6]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 3'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 3'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
        if( tscore[2] == 5'd0 && nextreqs[2] && (!busy || powner != 3'd2) )
          begin
            tscore_en[2]  = 1'b1;
            tscore_nxt[2] = nextqos[2];
          end
        if( tscore[3] == 5'd0 && nextreqs[3] && (!busy || powner != 3'd3) )
          begin
            tscore_en[3]  = 1'b1;
            tscore_nxt[3] = nextqos[3];
          end
        if( tscore[4] == 5'd0 && nextreqs[4] && (!busy || powner != 3'd4) )
          begin
            tscore_en[4]  = 1'b1;
            tscore_nxt[4] = nextqos[4];
          end
        if( tscore[5] == 5'd0 && nextreqs[5] && (!busy || powner != 3'd5) )
          begin
            tscore_en[5]  = 1'b1;
            tscore_nxt[5] = nextqos[5];
          end
        if( tscore[6] == 5'd0 && nextreqs[6] && (!busy || powner != 3'd6) )
          begin
            tscore_en[6]  = 1'b1;
            tscore_nxt[6] = nextqos[6];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign tmpMax1 = tscore_nxt[3]>tscore_nxt[2] ? tscore_nxt[3] : tscore_nxt[2];
assign tmpMax2 = tscore_nxt[5]>tscore_nxt[4] ? tscore_nxt[5] : tscore_nxt[4];
assign tmpMax3 = tscore_nxt[6]>tmpMax0 ? tscore_nxt[6] : tmpMax0;
assign tmpMax4 = tmpMax2>tmpMax1 ? tmpMax2 : tmpMax1;
assign tmpMax5 = tmpMax4>tmpMax3 ? tmpMax4 : tmpMax3;
assign maxScore_nxt = tmpMax5;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 7'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
  if( tscore[2]==maxScore )
    preqs[2] = prawreqs[2];
  if( tscore[3]==maxScore )
    preqs[3] = prawreqs[3];
  if( tscore[4]==maxScore )
    preqs[4] = prawreqs[4];
  if( tscore[5]==maxScore )
    preqs[5] = prawreqs[5];
  if( tscore[6]==maxScore )
    preqs[6] = prawreqs[6];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        3'd0: owner = (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 :  powner;
        3'd1: owner = (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 :  powner;
        3'd2: owner = (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 :  powner;
        3'd3: owner = (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 :  powner;
        3'd4: owner = (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 :  powner;
        3'd5: owner = (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 :  powner;
        3'd6: owner = (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    3'd0:
      begin
        int_flitdata = r0_t4_flitdata;
        int_sop      = r0_t4_sop;
        int_eop      = r0_t4_eop;
      end
    3'd1:
      begin
        int_flitdata = r0_t2_flitdata;
        int_sop      = r0_t2_sop;
        int_eop      = r0_t2_eop;
      end
    3'd2:
      begin
        int_flitdata = r0_t1_flitdata;
        int_sop      = r0_t1_sop;
        int_eop      = r0_t1_eop;
      end
    3'd3:
      begin
        int_flitdata = r0_t0_flitdata;
        int_sop      = r0_t0_sop;
        int_eop      = r0_t0_eop;
      end
    3'd4:
      begin
        int_flitdata = r0_t5_flitdata;
        int_sop      = r0_t5_sop;
        int_eop      = r0_t5_eop;
      end
    3'd5:
      begin
        int_flitdata = r0_t3_flitdata;
        int_sop      = r0_t3_sop;
        int_eop      = r0_t3_eop;
      end
    3'd6:
      begin
        int_flitdata = r0_t1000_flitdata;
        int_sop      = r0_t1000_sop;
        int_eop      = r0_t1000_eop;
      end
    default:
      begin
        int_flitdata = {34{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign r0_t4_i1_ready = int_ready && (owner == 3'd0);
assign r0_t2_i1_ready = int_ready && (owner == 3'd1);
assign r0_t1_i1_ready = int_ready && (owner == 3'd2);
assign r0_t0_i1_ready = int_ready && (owner == 3'd3);
assign r0_t5_i1_ready = int_ready && (owner == 3'd4);
assign r0_t3_i1_ready = int_ready && (owner == 3'd5);
assign r0_t1000_i1_ready = int_ready && (owner == 3'd6);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_r0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:34
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:34
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_RTR_INI0_r0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // r1_t4
  input  wire            r1_t4_sop,
  input  wire            r1_t4_eop,
  input  wire      [3:0] r1_t4_qos_nxt,
  input  wire      [3:0] r1_t4_qos,
  input  wire     [23:0] r1_t4_flitdata,
  input  wire            r1_t4_i1_activity,
  input  wire            r1_t4_i1_req_nxt,
  input  wire            r1_t4_i1_req,
  output logic           r1_t4_i1_ready,
  // r1_t2
  input  wire            r1_t2_sop,
  input  wire            r1_t2_eop,
  input  wire      [3:0] r1_t2_qos_nxt,
  input  wire      [3:0] r1_t2_qos,
  input  wire     [23:0] r1_t2_flitdata,
  input  wire            r1_t2_i1_activity,
  input  wire            r1_t2_i1_req_nxt,
  input  wire            r1_t2_i1_req,
  output logic           r1_t2_i1_ready,
  // r1_t1
  input  wire            r1_t1_sop,
  input  wire            r1_t1_eop,
  input  wire      [3:0] r1_t1_qos_nxt,
  input  wire      [3:0] r1_t1_qos,
  input  wire     [23:0] r1_t1_flitdata,
  input  wire            r1_t1_i1_activity,
  input  wire            r1_t1_i1_req_nxt,
  input  wire            r1_t1_i1_req,
  output logic           r1_t1_i1_ready,
  // r1_t0
  input  wire            r1_t0_sop,
  input  wire            r1_t0_eop,
  input  wire      [3:0] r1_t0_qos_nxt,
  input  wire      [3:0] r1_t0_qos,
  input  wire     [23:0] r1_t0_flitdata,
  input  wire            r1_t0_i1_activity,
  input  wire            r1_t0_i1_req_nxt,
  input  wire            r1_t0_i1_req,
  output logic           r1_t0_i1_ready,
  // r1_t5
  input  wire            r1_t5_sop,
  input  wire            r1_t5_eop,
  input  wire      [3:0] r1_t5_qos_nxt,
  input  wire      [3:0] r1_t5_qos,
  input  wire     [23:0] r1_t5_flitdata,
  input  wire            r1_t5_i1_activity,
  input  wire            r1_t5_i1_req_nxt,
  input  wire            r1_t5_i1_req,
  output logic           r1_t5_i1_ready,
  // r1_t3
  input  wire            r1_t3_sop,
  input  wire            r1_t3_eop,
  input  wire      [3:0] r1_t3_qos_nxt,
  input  wire      [3:0] r1_t3_qos,
  input  wire     [23:0] r1_t3_flitdata,
  input  wire            r1_t3_i1_activity,
  input  wire            r1_t3_i1_req_nxt,
  input  wire            r1_t3_i1_req,
  output logic           r1_t3_i1_ready,
  // r1_t1000
  input  wire            r1_t1000_sop,
  input  wire            r1_t1000_eop,
  input  wire      [3:0] r1_t1000_qos_nxt,
  input  wire      [3:0] r1_t1000_qos,
  input  wire     [23:0] r1_t1000_flitdata,
  input  wire            r1_t1000_i1_activity,
  input  wire            r1_t1000_i1_req_nxt,
  input  wire            r1_t1000_i1_req,
  output logic           r1_t1000_i1_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [23:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [23:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [6:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [6:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [6:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [6:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [6:0];
logic     [4:0] tscore_nxt [6:0];
logic     [6:0] tscore_en;
logic     [2:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [4:0] tmpMax1;
logic     [4:0] tmpMax2;
logic     [4:0] tmpMax3;
logic     [4:0] tmpMax4;
logic     [4:0] tmpMax5;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = r1_t4_i1_activity || r1_t4_i1_req || r1_t2_i1_activity || r1_t2_i1_req || r1_t1_i1_activity || r1_t1_i1_req || r1_t0_i1_activity || r1_t0_i1_req || r1_t5_i1_activity || r1_t5_i1_req || r1_t3_i1_activity || r1_t3_i1_req || r1_t1000_i1_activity || r1_t1000_i1_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_RTR_INI0_r1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
      tscore[2] <= #1ps 5'd0;
      tscore[3] <= #1ps 5'd0;
      tscore[4] <= #1ps 5'd0;
      tscore[5] <= #1ps 5'd0;
      tscore[6] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
      if (tscore_en[2])
        tscore[2] <= #1ps tscore_nxt[2];
      if (tscore_en[3])
        tscore[3] <= #1ps tscore_nxt[3];
      if (tscore_en[4])
        tscore[4] <= #1ps tscore_nxt[4];
      if (tscore_en[5])
        tscore[5] <= #1ps tscore_nxt[5];
      if (tscore_en[6])
        tscore[6] <= #1ps tscore_nxt[6];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 3'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = r1_t4_i1_req;
assign nextreqs[0] = r1_t4_i1_req_nxt;
assign nextqos[0] = r1_t4_qos_nxt + 4'd1;
assign prawreqs[1] = r1_t2_i1_req;
assign nextreqs[1] = r1_t2_i1_req_nxt;
assign nextqos[1] = r1_t2_qos_nxt + 4'd1;
assign prawreqs[2] = r1_t1_i1_req;
assign nextreqs[2] = r1_t1_i1_req_nxt;
assign nextqos[2] = r1_t1_qos_nxt + 4'd1;
assign prawreqs[3] = r1_t0_i1_req;
assign nextreqs[3] = r1_t0_i1_req_nxt;
assign nextqos[3] = r1_t0_qos_nxt + 4'd1;
assign prawreqs[4] = r1_t5_i1_req;
assign nextreqs[4] = r1_t5_i1_req_nxt;
assign nextqos[4] = r1_t5_qos_nxt + 4'd1;
assign prawreqs[5] = r1_t3_i1_req;
assign nextreqs[5] = r1_t3_i1_req_nxt;
assign nextqos[5] = r1_t3_qos_nxt + 4'd1;
assign prawreqs[6] = r1_t1000_i1_req;
assign nextreqs[6] = r1_t1000_i1_req_nxt;
assign nextqos[6] = r1_t1000_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_nxt[2] = tscore[2];
    tscore_nxt[3] = tscore[3];
    tscore_nxt[4] = tscore[4];
    tscore_nxt[5] = tscore[5];
    tscore_nxt[6] = tscore[6];
    tscore_en  = 7'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {7{1'b1}};
        if( owner==3'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==3'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
        if( owner==3'd2 || tscore[2] == 5'd0 )
          tscore_nxt[2] = nextreqs[2] ? nextqos[2] : 5'd0;
        else if( tscore[2]!=5'h1F )
          tscore_nxt[2] = tscore[2]+5'd1;
        if( owner==3'd3 || tscore[3] == 5'd0 )
          tscore_nxt[3] = nextreqs[3] ? nextqos[3] : 5'd0;
        else if( tscore[3]!=5'h1F )
          tscore_nxt[3] = tscore[3]+5'd1;
        if( owner==3'd4 || tscore[4] == 5'd0 )
          tscore_nxt[4] = nextreqs[4] ? nextqos[4] : 5'd0;
        else if( tscore[4]!=5'h1F )
          tscore_nxt[4] = tscore[4]+5'd1;
        if( owner==3'd5 || tscore[5] == 5'd0 )
          tscore_nxt[5] = nextreqs[5] ? nextqos[5] : 5'd0;
        else if( tscore[5]!=5'h1F )
          tscore_nxt[5] = tscore[5]+5'd1;
        if( owner==3'd6 || tscore[6] == 5'd0 )
          tscore_nxt[6] = nextreqs[6] ? nextqos[6] : 5'd0;
        else if( tscore[6]!=5'h1F )
          tscore_nxt[6] = tscore[6]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 3'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 3'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
        if( tscore[2] == 5'd0 && nextreqs[2] && (!busy || powner != 3'd2) )
          begin
            tscore_en[2]  = 1'b1;
            tscore_nxt[2] = nextqos[2];
          end
        if( tscore[3] == 5'd0 && nextreqs[3] && (!busy || powner != 3'd3) )
          begin
            tscore_en[3]  = 1'b1;
            tscore_nxt[3] = nextqos[3];
          end
        if( tscore[4] == 5'd0 && nextreqs[4] && (!busy || powner != 3'd4) )
          begin
            tscore_en[4]  = 1'b1;
            tscore_nxt[4] = nextqos[4];
          end
        if( tscore[5] == 5'd0 && nextreqs[5] && (!busy || powner != 3'd5) )
          begin
            tscore_en[5]  = 1'b1;
            tscore_nxt[5] = nextqos[5];
          end
        if( tscore[6] == 5'd0 && nextreqs[6] && (!busy || powner != 3'd6) )
          begin
            tscore_en[6]  = 1'b1;
            tscore_nxt[6] = nextqos[6];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign tmpMax1 = tscore_nxt[3]>tscore_nxt[2] ? tscore_nxt[3] : tscore_nxt[2];
assign tmpMax2 = tscore_nxt[5]>tscore_nxt[4] ? tscore_nxt[5] : tscore_nxt[4];
assign tmpMax3 = tscore_nxt[6]>tmpMax0 ? tscore_nxt[6] : tmpMax0;
assign tmpMax4 = tmpMax2>tmpMax1 ? tmpMax2 : tmpMax1;
assign tmpMax5 = tmpMax4>tmpMax3 ? tmpMax4 : tmpMax3;
assign maxScore_nxt = tmpMax5;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 7'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
  if( tscore[2]==maxScore )
    preqs[2] = prawreqs[2];
  if( tscore[3]==maxScore )
    preqs[3] = prawreqs[3];
  if( tscore[4]==maxScore )
    preqs[4] = prawreqs[4];
  if( tscore[5]==maxScore )
    preqs[5] = prawreqs[5];
  if( tscore[6]==maxScore )
    preqs[6] = prawreqs[6];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        3'd0: owner = (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 :  powner;
        3'd1: owner = (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 :  powner;
        3'd2: owner = (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 :  powner;
        3'd3: owner = (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 :  powner;
        3'd4: owner = (preqs[5]) ? 3'd5 : (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 :  powner;
        3'd5: owner = (preqs[6]) ? 3'd6 : (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 :  powner;
        3'd6: owner = (preqs[0]) ? 3'd0 : (preqs[1]) ? 3'd1 : (preqs[2]) ? 3'd2 : (preqs[3]) ? 3'd3 : (preqs[4]) ? 3'd4 : (preqs[5]) ? 3'd5 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    3'd0:
      begin
        int_flitdata = r1_t4_flitdata;
        int_sop      = r1_t4_sop;
        int_eop      = r1_t4_eop;
      end
    3'd1:
      begin
        int_flitdata = r1_t2_flitdata;
        int_sop      = r1_t2_sop;
        int_eop      = r1_t2_eop;
      end
    3'd2:
      begin
        int_flitdata = r1_t1_flitdata;
        int_sop      = r1_t1_sop;
        int_eop      = r1_t1_eop;
      end
    3'd3:
      begin
        int_flitdata = r1_t0_flitdata;
        int_sop      = r1_t0_sop;
        int_eop      = r1_t0_eop;
      end
    3'd4:
      begin
        int_flitdata = r1_t5_flitdata;
        int_sop      = r1_t5_sop;
        int_eop      = r1_t5_eop;
      end
    3'd5:
      begin
        int_flitdata = r1_t3_flitdata;
        int_sop      = r1_t3_sop;
        int_eop      = r1_t3_eop;
      end
    3'd6:
      begin
        int_flitdata = r1_t1000_flitdata;
        int_sop      = r1_t1000_sop;
        int_eop      = r1_t1000_eop;
      end
    default:
      begin
        int_flitdata = {24{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign r1_t4_i1_ready = int_ready && (owner == 3'd0);
assign r1_t2_i1_ready = int_ready && (owner == 3'd1);
assign r1_t1_i1_ready = int_ready && (owner == 3'd2);
assign r1_t0_i1_ready = int_ready && (owner == 3'd3);
assign r1_t5_i1_ready = int_ready && (owner == 3'd4);
assign r1_t3_i1_ready = int_ready && (owner == 3'd5);
assign r1_t1000_i1_ready = int_ready && (owner == 3'd6);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_RTR_INI0_r1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:24
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:24
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_RTR_INI0_r1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_RTR_INI0_r1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f0_i0
  input  wire            f0_i0_sop,
  input  wire            f0_i0_eop,
  input  wire      [3:0] f0_i0_qos_nxt,
  input  wire      [3:0] f0_i0_qos,
  input  wire     [35:0] f0_i0_flitdata,
  input  wire            f0_i0_t0_activity,
  input  wire            f0_i0_t0_req_nxt,
  input  wire            f0_i0_t0_req,
  output logic           f0_i0_t0_ready,
  // f0_i1
  input  wire            f0_i1_sop,
  input  wire            f0_i1_eop,
  input  wire      [3:0] f0_i1_qos_nxt,
  input  wire      [3:0] f0_i1_qos,
  input  wire     [35:0] f0_i1_flitdata,
  input  wire            f0_i1_t0_activity,
  input  wire            f0_i1_t0_req_nxt,
  input  wire            f0_i1_t0_req,
  output logic           f0_i1_t0_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [35:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [35:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f0_i0_t0_activity || f0_i0_t0_req || f0_i1_t0_activity || f0_i1_t0_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f0_i0_t0_req;
assign nextreqs[0] = f0_i0_t0_req_nxt;
assign nextqos[0] = f0_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f0_i1_t0_req;
assign nextreqs[1] = f0_i1_t0_req_nxt;
assign nextqos[1] = f0_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f0_i0_flitdata;
        int_sop      = f0_i0_sop;
        int_eop      = f0_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f0_i1_flitdata;
        int_sop      = f0_i1_sop;
        int_eop      = f0_i1_eop;
      end
    default:
      begin
        int_flitdata = {36{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f0_i0_t0_ready = int_ready && (owner == 1'd0);
assign f0_i1_t0_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:36
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:36
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f1_i0
  input  wire            f1_i0_sop,
  input  wire            f1_i0_eop,
  input  wire      [3:0] f1_i0_qos_nxt,
  input  wire      [3:0] f1_i0_qos,
  input  wire     [59:0] f1_i0_flitdata,
  input  wire            f1_i0_t0_activity,
  input  wire            f1_i0_t0_req_nxt,
  input  wire            f1_i0_t0_req,
  output logic           f1_i0_t0_ready,
  // f1_i1
  input  wire            f1_i1_sop,
  input  wire            f1_i1_eop,
  input  wire      [3:0] f1_i1_qos_nxt,
  input  wire      [3:0] f1_i1_qos,
  input  wire     [59:0] f1_i1_flitdata,
  input  wire            f1_i1_t0_activity,
  input  wire            f1_i1_t0_req_nxt,
  input  wire            f1_i1_t0_req,
  output logic           f1_i1_t0_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [59:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [59:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f1_i0_t0_activity || f1_i0_t0_req || f1_i1_t0_activity || f1_i1_t0_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f1_i0_t0_req;
assign nextreqs[0] = f1_i0_t0_req_nxt;
assign nextqos[0] = f1_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f1_i1_t0_req;
assign nextreqs[1] = f1_i1_t0_req_nxt;
assign nextqos[1] = f1_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f1_i0_flitdata;
        int_sop      = f1_i0_sop;
        int_eop      = f1_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f1_i1_flitdata;
        int_sop      = f1_i1_sop;
        int_eop      = f1_i1_eop;
      end
    default:
      begin
        int_flitdata = {60{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f1_i0_t0_ready = int_ready && (owner == 1'd0);
assign f1_i1_t0_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:60
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:60
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_f1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [33:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r0_t0
  output logic           r0_t0_sop,
  output logic           r0_t0_eop,
  output logic     [3:0] r0_t0_qos_nxt,
  output logic     [3:0] r0_t0_qos,
  output logic    [33:0] r0_t0_flitdata,
  output logic           r0_t0_i0_activity,
  output logic           r0_t0_i0_req_nxt,
  output logic           r0_t0_i0_req,
  input  wire            r0_t0_i0_ready,
  output logic           r0_t0_i1_activity,
  output logic           r0_t0_i1_req_nxt,
  output logic           r0_t0_i1_req,
  input  wire            r0_t0_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [33:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [33:0] intp_flitdata;
logic    [33:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:34
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:34
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r0_t0_i0_req = tgtReq[1];
assign tgtXfer[1] = r0_t0_i0_req && r0_t0_i0_ready;
assign r0_t0_i0_activity = tgtAct[1];
assign r0_t0_i0_req_nxt = tgtReqNxt[1];
assign r0_t0_i1_req = tgtReq[0];
assign tgtXfer[0] = r0_t0_i1_req && r0_t0_i1_ready;
assign r0_t0_i1_activity = tgtAct[0];
assign r0_t0_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:34
  .intp_flitdata(intp_flitdata),                                                // o:34
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:34
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r0_t0_sop = intp_sop;
assign r0_t0_eop = intp_eop;
assign r0_t0_qos = intp_qos;
assign r0_t0_flitdata = intp_flitdata;
assign r0_t0_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [33:0] int_flitdata,
  output logic    [33:0] intp_flitdata,
  output logic    [33:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [40:0] wdata;
logic    [40:0] rdata;
logic    [40:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [40:0] fifodata [1:0];
logic    [40:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[35:2] = int_flitdata;
assign intp_flitdata = rdata[35:2];
assign intp_flitdata_nxt = rdata_nxt[35:2];
assign wdata[39:36] = int_qos;
assign intp_qos = rdata[39:36];
assign intp_qos_nxt = rdata_nxt[39:36];
assign wdata[40:40] = int_dstIdx;
assign intp_dstIdx = rdata[40:40];
assign intp_dstIdx_nxt = rdata_nxt[40:40];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {41{1'b0}};
      fifodata[1] <= #1ps {41{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {41{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [23:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r1_t0
  output logic           r1_t0_sop,
  output logic           r1_t0_eop,
  output logic     [3:0] r1_t0_qos_nxt,
  output logic     [3:0] r1_t0_qos,
  output logic    [23:0] r1_t0_flitdata,
  output logic           r1_t0_i0_activity,
  output logic           r1_t0_i0_req_nxt,
  output logic           r1_t0_i0_req,
  input  wire            r1_t0_i0_ready,
  output logic           r1_t0_i1_activity,
  output logic           r1_t0_i1_req_nxt,
  output logic           r1_t0_i1_req,
  input  wire            r1_t0_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [23:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [23:0] intp_flitdata;
logic    [23:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:24
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:24
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r1_t0_i0_req = tgtReq[1];
assign tgtXfer[1] = r1_t0_i0_req && r1_t0_i0_ready;
assign r1_t0_i0_activity = tgtAct[1];
assign r1_t0_i0_req_nxt = tgtReqNxt[1];
assign r1_t0_i1_req = tgtReq[0];
assign tgtXfer[0] = r1_t0_i1_req && r1_t0_i1_ready;
assign r1_t0_i1_activity = tgtAct[0];
assign r1_t0_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:24
  .intp_flitdata(intp_flitdata),                                                // o:24
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:24
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r1_t0_sop = intp_sop;
assign r1_t0_eop = intp_eop;
assign r1_t0_qos = intp_qos;
assign r1_t0_flitdata = intp_flitdata;
assign r1_t0_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [23:0] int_flitdata,
  output logic    [23:0] intp_flitdata,
  output logic    [23:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [30:0] wdata;
logic    [30:0] rdata;
logic    [30:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [30:0] fifodata [1:0];
logic    [30:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[25:2] = int_flitdata;
assign intp_flitdata = rdata[25:2];
assign intp_flitdata_nxt = rdata_nxt[25:2];
assign wdata[29:26] = int_qos;
assign intp_qos = rdata[29:26];
assign intp_qos_nxt = rdata_nxt[29:26];
assign wdata[30:30] = int_dstIdx;
assign intp_dstIdx = rdata[30:30];
assign intp_dstIdx_nxt = rdata_nxt[30:30];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps 31'd0;
      fifodata[1] <= #1ps 31'd0;
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {31{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_cmn_TEA_r1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f0_i0
  input  wire            f0_i0_sop,
  input  wire            f0_i0_eop,
  input  wire      [3:0] f0_i0_qos_nxt,
  input  wire      [3:0] f0_i0_qos,
  input  wire     [35:0] f0_i0_flitdata,
  input  wire            f0_i0_t1_activity,
  input  wire            f0_i0_t1_req_nxt,
  input  wire            f0_i0_t1_req,
  output logic           f0_i0_t1_ready,
  // f0_i1
  input  wire            f0_i1_sop,
  input  wire            f0_i1_eop,
  input  wire      [3:0] f0_i1_qos_nxt,
  input  wire      [3:0] f0_i1_qos,
  input  wire     [35:0] f0_i1_flitdata,
  input  wire            f0_i1_t1_activity,
  input  wire            f0_i1_t1_req_nxt,
  input  wire            f0_i1_t1_req,
  output logic           f0_i1_t1_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [35:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [35:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f0_i0_t1_activity || f0_i0_t1_req || f0_i1_t1_activity || f0_i1_t1_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f0_i0_t1_req;
assign nextreqs[0] = f0_i0_t1_req_nxt;
assign nextqos[0] = f0_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f0_i1_t1_req;
assign nextreqs[1] = f0_i1_t1_req_nxt;
assign nextqos[1] = f0_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f0_i0_flitdata;
        int_sop      = f0_i0_sop;
        int_eop      = f0_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f0_i1_flitdata;
        int_sop      = f0_i1_sop;
        int_eop      = f0_i1_eop;
      end
    default:
      begin
        int_flitdata = {36{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f0_i0_t1_ready = int_ready && (owner == 1'd0);
assign f0_i1_t1_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:36
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:36
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f1_i0
  input  wire            f1_i0_sop,
  input  wire            f1_i0_eop,
  input  wire      [3:0] f1_i0_qos_nxt,
  input  wire      [3:0] f1_i0_qos,
  input  wire     [59:0] f1_i0_flitdata,
  input  wire            f1_i0_t1_activity,
  input  wire            f1_i0_t1_req_nxt,
  input  wire            f1_i0_t1_req,
  output logic           f1_i0_t1_ready,
  // f1_i1
  input  wire            f1_i1_sop,
  input  wire            f1_i1_eop,
  input  wire      [3:0] f1_i1_qos_nxt,
  input  wire      [3:0] f1_i1_qos,
  input  wire     [59:0] f1_i1_flitdata,
  input  wire            f1_i1_t1_activity,
  input  wire            f1_i1_t1_req_nxt,
  input  wire            f1_i1_t1_req,
  output logic           f1_i1_t1_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [59:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [59:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f1_i0_t1_activity || f1_i0_t1_req || f1_i1_t1_activity || f1_i1_t1_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f1_i0_t1_req;
assign nextreqs[0] = f1_i0_t1_req_nxt;
assign nextqos[0] = f1_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f1_i1_t1_req;
assign nextreqs[1] = f1_i1_t1_req_nxt;
assign nextqos[1] = f1_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f1_i0_flitdata;
        int_sop      = f1_i0_sop;
        int_eop      = f1_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f1_i1_flitdata;
        int_sop      = f1_i1_sop;
        int_eop      = f1_i1_eop;
      end
    default:
      begin
        int_flitdata = {60{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f1_i0_t1_ready = int_ready && (owner == 1'd0);
assign f1_i1_t1_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:60
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:60
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_f1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [33:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r0_t1
  output logic           r0_t1_sop,
  output logic           r0_t1_eop,
  output logic     [3:0] r0_t1_qos_nxt,
  output logic     [3:0] r0_t1_qos,
  output logic    [33:0] r0_t1_flitdata,
  output logic           r0_t1_i0_activity,
  output logic           r0_t1_i0_req_nxt,
  output logic           r0_t1_i0_req,
  input  wire            r0_t1_i0_ready,
  output logic           r0_t1_i1_activity,
  output logic           r0_t1_i1_req_nxt,
  output logic           r0_t1_i1_req,
  input  wire            r0_t1_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [33:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [33:0] intp_flitdata;
logic    [33:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:34
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:34
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r0_t1_i0_req = tgtReq[1];
assign tgtXfer[1] = r0_t1_i0_req && r0_t1_i0_ready;
assign r0_t1_i0_activity = tgtAct[1];
assign r0_t1_i0_req_nxt = tgtReqNxt[1];
assign r0_t1_i1_req = tgtReq[0];
assign tgtXfer[0] = r0_t1_i1_req && r0_t1_i1_ready;
assign r0_t1_i1_activity = tgtAct[0];
assign r0_t1_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:34
  .intp_flitdata(intp_flitdata),                                                // o:34
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:34
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r0_t1_sop = intp_sop;
assign r0_t1_eop = intp_eop;
assign r0_t1_qos = intp_qos;
assign r0_t1_flitdata = intp_flitdata;
assign r0_t1_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [33:0] int_flitdata,
  output logic    [33:0] intp_flitdata,
  output logic    [33:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [40:0] wdata;
logic    [40:0] rdata;
logic    [40:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [40:0] fifodata [1:0];
logic    [40:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[35:2] = int_flitdata;
assign intp_flitdata = rdata[35:2];
assign intp_flitdata_nxt = rdata_nxt[35:2];
assign wdata[39:36] = int_qos;
assign intp_qos = rdata[39:36];
assign intp_qos_nxt = rdata_nxt[39:36];
assign wdata[40:40] = int_dstIdx;
assign intp_dstIdx = rdata[40:40];
assign intp_dstIdx_nxt = rdata_nxt[40:40];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {41{1'b0}};
      fifodata[1] <= #1ps {41{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {41{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [23:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r1_t1
  output logic           r1_t1_sop,
  output logic           r1_t1_eop,
  output logic     [3:0] r1_t1_qos_nxt,
  output logic     [3:0] r1_t1_qos,
  output logic    [23:0] r1_t1_flitdata,
  output logic           r1_t1_i0_activity,
  output logic           r1_t1_i0_req_nxt,
  output logic           r1_t1_i0_req,
  input  wire            r1_t1_i0_ready,
  output logic           r1_t1_i1_activity,
  output logic           r1_t1_i1_req_nxt,
  output logic           r1_t1_i1_req,
  input  wire            r1_t1_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [23:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [23:0] intp_flitdata;
logic    [23:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:24
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:24
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r1_t1_i0_req = tgtReq[1];
assign tgtXfer[1] = r1_t1_i0_req && r1_t1_i0_ready;
assign r1_t1_i0_activity = tgtAct[1];
assign r1_t1_i0_req_nxt = tgtReqNxt[1];
assign r1_t1_i1_req = tgtReq[0];
assign tgtXfer[0] = r1_t1_i1_req && r1_t1_i1_ready;
assign r1_t1_i1_activity = tgtAct[0];
assign r1_t1_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:24
  .intp_flitdata(intp_flitdata),                                                // o:24
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:24
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r1_t1_sop = intp_sop;
assign r1_t1_eop = intp_eop;
assign r1_t1_qos = intp_qos;
assign r1_t1_flitdata = intp_flitdata;
assign r1_t1_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [23:0] int_flitdata,
  output logic    [23:0] intp_flitdata,
  output logic    [23:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [30:0] wdata;
logic    [30:0] rdata;
logic    [30:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [30:0] fifodata [1:0];
logic    [30:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[25:2] = int_flitdata;
assign intp_flitdata = rdata[25:2];
assign intp_flitdata_nxt = rdata_nxt[25:2];
assign wdata[29:26] = int_qos;
assign intp_qos = rdata[29:26];
assign intp_qos_nxt = rdata_nxt[29:26];
assign wdata[30:30] = int_dstIdx;
assign intp_dstIdx = rdata[30:30];
assign intp_dstIdx_nxt = rdata_nxt[30:30];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps 31'd0;
      fifodata[1] <= #1ps 31'd0;
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {31{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_tc_reg_TEA_r1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f0_i0
  input  wire            f0_i0_sop,
  input  wire            f0_i0_eop,
  input  wire      [3:0] f0_i0_qos_nxt,
  input  wire      [3:0] f0_i0_qos,
  input  wire     [35:0] f0_i0_flitdata,
  input  wire            f0_i0_t2_activity,
  input  wire            f0_i0_t2_req_nxt,
  input  wire            f0_i0_t2_req,
  output logic           f0_i0_t2_ready,
  // f0_i1
  input  wire            f0_i1_sop,
  input  wire            f0_i1_eop,
  input  wire      [3:0] f0_i1_qos_nxt,
  input  wire      [3:0] f0_i1_qos,
  input  wire     [35:0] f0_i1_flitdata,
  input  wire            f0_i1_t2_activity,
  input  wire            f0_i1_t2_req_nxt,
  input  wire            f0_i1_t2_req,
  output logic           f0_i1_t2_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [35:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [35:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f0_i0_t2_activity || f0_i0_t2_req || f0_i1_t2_activity || f0_i1_t2_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f0_i0_t2_req;
assign nextreqs[0] = f0_i0_t2_req_nxt;
assign nextqos[0] = f0_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f0_i1_t2_req;
assign nextreqs[1] = f0_i1_t2_req_nxt;
assign nextqos[1] = f0_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f0_i0_flitdata;
        int_sop      = f0_i0_sop;
        int_eop      = f0_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f0_i1_flitdata;
        int_sop      = f0_i1_sop;
        int_eop      = f0_i1_eop;
      end
    default:
      begin
        int_flitdata = {36{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f0_i0_t2_ready = int_ready && (owner == 1'd0);
assign f0_i1_t2_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:36
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:36
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f1_i0
  input  wire            f1_i0_sop,
  input  wire            f1_i0_eop,
  input  wire      [3:0] f1_i0_qos_nxt,
  input  wire      [3:0] f1_i0_qos,
  input  wire     [59:0] f1_i0_flitdata,
  input  wire            f1_i0_t2_activity,
  input  wire            f1_i0_t2_req_nxt,
  input  wire            f1_i0_t2_req,
  output logic           f1_i0_t2_ready,
  // f1_i1
  input  wire            f1_i1_sop,
  input  wire            f1_i1_eop,
  input  wire      [3:0] f1_i1_qos_nxt,
  input  wire      [3:0] f1_i1_qos,
  input  wire     [59:0] f1_i1_flitdata,
  input  wire            f1_i1_t2_activity,
  input  wire            f1_i1_t2_req_nxt,
  input  wire            f1_i1_t2_req,
  output logic           f1_i1_t2_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [59:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [59:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f1_i0_t2_activity || f1_i0_t2_req || f1_i1_t2_activity || f1_i1_t2_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f1_i0_t2_req;
assign nextreqs[0] = f1_i0_t2_req_nxt;
assign nextqos[0] = f1_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f1_i1_t2_req;
assign nextreqs[1] = f1_i1_t2_req_nxt;
assign nextqos[1] = f1_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f1_i0_flitdata;
        int_sop      = f1_i0_sop;
        int_eop      = f1_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f1_i1_flitdata;
        int_sop      = f1_i1_sop;
        int_eop      = f1_i1_eop;
      end
    default:
      begin
        int_flitdata = {60{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f1_i0_t2_ready = int_ready && (owner == 1'd0);
assign f1_i1_t2_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:60
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:60
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_f1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [33:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r0_t2
  output logic           r0_t2_sop,
  output logic           r0_t2_eop,
  output logic     [3:0] r0_t2_qos_nxt,
  output logic     [3:0] r0_t2_qos,
  output logic    [33:0] r0_t2_flitdata,
  output logic           r0_t2_i0_activity,
  output logic           r0_t2_i0_req_nxt,
  output logic           r0_t2_i0_req,
  input  wire            r0_t2_i0_ready,
  output logic           r0_t2_i1_activity,
  output logic           r0_t2_i1_req_nxt,
  output logic           r0_t2_i1_req,
  input  wire            r0_t2_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [33:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [33:0] intp_flitdata;
logic    [33:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:34
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:34
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r0_t2_i0_req = tgtReq[1];
assign tgtXfer[1] = r0_t2_i0_req && r0_t2_i0_ready;
assign r0_t2_i0_activity = tgtAct[1];
assign r0_t2_i0_req_nxt = tgtReqNxt[1];
assign r0_t2_i1_req = tgtReq[0];
assign tgtXfer[0] = r0_t2_i1_req && r0_t2_i1_ready;
assign r0_t2_i1_activity = tgtAct[0];
assign r0_t2_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:34
  .intp_flitdata(intp_flitdata),                                                // o:34
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:34
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r0_t2_sop = intp_sop;
assign r0_t2_eop = intp_eop;
assign r0_t2_qos = intp_qos;
assign r0_t2_flitdata = intp_flitdata;
assign r0_t2_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [33:0] int_flitdata,
  output logic    [33:0] intp_flitdata,
  output logic    [33:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [40:0] wdata;
logic    [40:0] rdata;
logic    [40:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [40:0] fifodata [1:0];
logic    [40:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[35:2] = int_flitdata;
assign intp_flitdata = rdata[35:2];
assign intp_flitdata_nxt = rdata_nxt[35:2];
assign wdata[39:36] = int_qos;
assign intp_qos = rdata[39:36];
assign intp_qos_nxt = rdata_nxt[39:36];
assign wdata[40:40] = int_dstIdx;
assign intp_dstIdx = rdata[40:40];
assign intp_dstIdx_nxt = rdata_nxt[40:40];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {41{1'b0}};
      fifodata[1] <= #1ps {41{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {41{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [23:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r1_t2
  output logic           r1_t2_sop,
  output logic           r1_t2_eop,
  output logic     [3:0] r1_t2_qos_nxt,
  output logic     [3:0] r1_t2_qos,
  output logic    [23:0] r1_t2_flitdata,
  output logic           r1_t2_i0_activity,
  output logic           r1_t2_i0_req_nxt,
  output logic           r1_t2_i0_req,
  input  wire            r1_t2_i0_ready,
  output logic           r1_t2_i1_activity,
  output logic           r1_t2_i1_req_nxt,
  output logic           r1_t2_i1_req,
  input  wire            r1_t2_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [23:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [23:0] intp_flitdata;
logic    [23:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:24
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:24
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r1_t2_i0_req = tgtReq[1];
assign tgtXfer[1] = r1_t2_i0_req && r1_t2_i0_ready;
assign r1_t2_i0_activity = tgtAct[1];
assign r1_t2_i0_req_nxt = tgtReqNxt[1];
assign r1_t2_i1_req = tgtReq[0];
assign tgtXfer[0] = r1_t2_i1_req && r1_t2_i1_ready;
assign r1_t2_i1_activity = tgtAct[0];
assign r1_t2_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:24
  .intp_flitdata(intp_flitdata),                                                // o:24
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:24
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r1_t2_sop = intp_sop;
assign r1_t2_eop = intp_eop;
assign r1_t2_qos = intp_qos;
assign r1_t2_flitdata = intp_flitdata;
assign r1_t2_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [23:0] int_flitdata,
  output logic    [23:0] intp_flitdata,
  output logic    [23:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [30:0] wdata;
logic    [30:0] rdata;
logic    [30:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [30:0] fifodata [1:0];
logic    [30:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[25:2] = int_flitdata;
assign intp_flitdata = rdata[25:2];
assign intp_flitdata_nxt = rdata_nxt[25:2];
assign wdata[29:26] = int_qos;
assign intp_qos = rdata[29:26];
assign intp_qos_nxt = rdata_nxt[29:26];
assign wdata[30:30] = int_dstIdx;
assign intp_dstIdx = rdata[30:30];
assign intp_dstIdx_nxt = rdata_nxt[30:30];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps 31'd0;
      fifodata[1] <= #1ps 31'd0;
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {31{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb_sub_sys_TEA_r1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f0_i0
  input  wire            f0_i0_sop,
  input  wire            f0_i0_eop,
  input  wire      [3:0] f0_i0_qos_nxt,
  input  wire      [3:0] f0_i0_qos,
  input  wire     [35:0] f0_i0_flitdata,
  input  wire            f0_i0_t3_activity,
  input  wire            f0_i0_t3_req_nxt,
  input  wire            f0_i0_t3_req,
  output logic           f0_i0_t3_ready,
  // f0_i1
  input  wire            f0_i1_sop,
  input  wire            f0_i1_eop,
  input  wire      [3:0] f0_i1_qos_nxt,
  input  wire      [3:0] f0_i1_qos,
  input  wire     [35:0] f0_i1_flitdata,
  input  wire            f0_i1_t3_activity,
  input  wire            f0_i1_t3_req_nxt,
  input  wire            f0_i1_t3_req,
  output logic           f0_i1_t3_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [35:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [35:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f0_i0_t3_activity || f0_i0_t3_req || f0_i1_t3_activity || f0_i1_t3_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f0_i0_t3_req;
assign nextreqs[0] = f0_i0_t3_req_nxt;
assign nextqos[0] = f0_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f0_i1_t3_req;
assign nextreqs[1] = f0_i1_t3_req_nxt;
assign nextqos[1] = f0_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f0_i0_flitdata;
        int_sop      = f0_i0_sop;
        int_eop      = f0_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f0_i1_flitdata;
        int_sop      = f0_i1_sop;
        int_eop      = f0_i1_eop;
      end
    default:
      begin
        int_flitdata = {36{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f0_i0_t3_ready = int_ready && (owner == 1'd0);
assign f0_i1_t3_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:36
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:36
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f1_i0
  input  wire            f1_i0_sop,
  input  wire            f1_i0_eop,
  input  wire      [3:0] f1_i0_qos_nxt,
  input  wire      [3:0] f1_i0_qos,
  input  wire     [59:0] f1_i0_flitdata,
  input  wire            f1_i0_t3_activity,
  input  wire            f1_i0_t3_req_nxt,
  input  wire            f1_i0_t3_req,
  output logic           f1_i0_t3_ready,
  // f1_i1
  input  wire            f1_i1_sop,
  input  wire            f1_i1_eop,
  input  wire      [3:0] f1_i1_qos_nxt,
  input  wire      [3:0] f1_i1_qos,
  input  wire     [59:0] f1_i1_flitdata,
  input  wire            f1_i1_t3_activity,
  input  wire            f1_i1_t3_req_nxt,
  input  wire            f1_i1_t3_req,
  output logic           f1_i1_t3_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [59:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [59:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f1_i0_t3_activity || f1_i0_t3_req || f1_i1_t3_activity || f1_i1_t3_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f1_i0_t3_req;
assign nextreqs[0] = f1_i0_t3_req_nxt;
assign nextqos[0] = f1_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f1_i1_t3_req;
assign nextreqs[1] = f1_i1_t3_req_nxt;
assign nextqos[1] = f1_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f1_i0_flitdata;
        int_sop      = f1_i0_sop;
        int_eop      = f1_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f1_i1_flitdata;
        int_sop      = f1_i1_sop;
        int_eop      = f1_i1_eop;
      end
    default:
      begin
        int_flitdata = {60{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f1_i0_t3_ready = int_ready && (owner == 1'd0);
assign f1_i1_t3_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:60
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:60
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_f1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [33:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r0_t3
  output logic           r0_t3_sop,
  output logic           r0_t3_eop,
  output logic     [3:0] r0_t3_qos_nxt,
  output logic     [3:0] r0_t3_qos,
  output logic    [33:0] r0_t3_flitdata,
  output logic           r0_t3_i0_activity,
  output logic           r0_t3_i0_req_nxt,
  output logic           r0_t3_i0_req,
  input  wire            r0_t3_i0_ready,
  output logic           r0_t3_i1_activity,
  output logic           r0_t3_i1_req_nxt,
  output logic           r0_t3_i1_req,
  input  wire            r0_t3_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [33:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [33:0] intp_flitdata;
logic    [33:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:34
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:34
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r0_t3_i0_req = tgtReq[1];
assign tgtXfer[1] = r0_t3_i0_req && r0_t3_i0_ready;
assign r0_t3_i0_activity = tgtAct[1];
assign r0_t3_i0_req_nxt = tgtReqNxt[1];
assign r0_t3_i1_req = tgtReq[0];
assign tgtXfer[0] = r0_t3_i1_req && r0_t3_i1_ready;
assign r0_t3_i1_activity = tgtAct[0];
assign r0_t3_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:34
  .intp_flitdata(intp_flitdata),                                                // o:34
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:34
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r0_t3_sop = intp_sop;
assign r0_t3_eop = intp_eop;
assign r0_t3_qos = intp_qos;
assign r0_t3_flitdata = intp_flitdata;
assign r0_t3_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [33:0] int_flitdata,
  output logic    [33:0] intp_flitdata,
  output logic    [33:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [40:0] wdata;
logic    [40:0] rdata;
logic    [40:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [40:0] fifodata [1:0];
logic    [40:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[35:2] = int_flitdata;
assign intp_flitdata = rdata[35:2];
assign intp_flitdata_nxt = rdata_nxt[35:2];
assign wdata[39:36] = int_qos;
assign intp_qos = rdata[39:36];
assign intp_qos_nxt = rdata_nxt[39:36];
assign wdata[40:40] = int_dstIdx;
assign intp_dstIdx = rdata[40:40];
assign intp_dstIdx_nxt = rdata_nxt[40:40];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {41{1'b0}};
      fifodata[1] <= #1ps {41{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {41{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [23:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r1_t3
  output logic           r1_t3_sop,
  output logic           r1_t3_eop,
  output logic     [3:0] r1_t3_qos_nxt,
  output logic     [3:0] r1_t3_qos,
  output logic    [23:0] r1_t3_flitdata,
  output logic           r1_t3_i0_activity,
  output logic           r1_t3_i0_req_nxt,
  output logic           r1_t3_i0_req,
  input  wire            r1_t3_i0_ready,
  output logic           r1_t3_i1_activity,
  output logic           r1_t3_i1_req_nxt,
  output logic           r1_t3_i1_req,
  input  wire            r1_t3_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [23:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [23:0] intp_flitdata;
logic    [23:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:24
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:24
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r1_t3_i0_req = tgtReq[1];
assign tgtXfer[1] = r1_t3_i0_req && r1_t3_i0_ready;
assign r1_t3_i0_activity = tgtAct[1];
assign r1_t3_i0_req_nxt = tgtReqNxt[1];
assign r1_t3_i1_req = tgtReq[0];
assign tgtXfer[0] = r1_t3_i1_req && r1_t3_i1_ready;
assign r1_t3_i1_activity = tgtAct[0];
assign r1_t3_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:24
  .intp_flitdata(intp_flitdata),                                                // o:24
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:24
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r1_t3_sop = intp_sop;
assign r1_t3_eop = intp_eop;
assign r1_t3_qos = intp_qos;
assign r1_t3_flitdata = intp_flitdata;
assign r1_t3_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [23:0] int_flitdata,
  output logic    [23:0] intp_flitdata,
  output logic    [23:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [30:0] wdata;
logic    [30:0] rdata;
logic    [30:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [30:0] fifodata [1:0];
logic    [30:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[25:2] = int_flitdata;
assign intp_flitdata = rdata[25:2];
assign intp_flitdata_nxt = rdata_nxt[25:2];
assign wdata[29:26] = int_qos;
assign intp_qos = rdata[29:26];
assign intp_qos_nxt = rdata_nxt[29:26];
assign wdata[30:30] = int_dstIdx;
assign intp_dstIdx = rdata[30:30];
assign intp_dstIdx_nxt = rdata_nxt[30:30];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps 31'd0;
      fifodata[1] <= #1ps 31'd0;
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {31{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_sub_sys_TEA_r1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f0_i0
  input  wire            f0_i0_sop,
  input  wire            f0_i0_eop,
  input  wire      [3:0] f0_i0_qos_nxt,
  input  wire      [3:0] f0_i0_qos,
  input  wire     [35:0] f0_i0_flitdata,
  input  wire            f0_i0_t4_activity,
  input  wire            f0_i0_t4_req_nxt,
  input  wire            f0_i0_t4_req,
  output logic           f0_i0_t4_ready,
  // f0_i1
  input  wire            f0_i1_sop,
  input  wire            f0_i1_eop,
  input  wire      [3:0] f0_i1_qos_nxt,
  input  wire      [3:0] f0_i1_qos,
  input  wire     [35:0] f0_i1_flitdata,
  input  wire            f0_i1_t4_activity,
  input  wire            f0_i1_t4_req_nxt,
  input  wire            f0_i1_t4_req,
  output logic           f0_i1_t4_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [35:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [35:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f0_i0_t4_activity || f0_i0_t4_req || f0_i1_t4_activity || f0_i1_t4_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f0_i0_t4_req;
assign nextreqs[0] = f0_i0_t4_req_nxt;
assign nextqos[0] = f0_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f0_i1_t4_req;
assign nextreqs[1] = f0_i1_t4_req_nxt;
assign nextqos[1] = f0_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f0_i0_flitdata;
        int_sop      = f0_i0_sop;
        int_eop      = f0_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f0_i1_flitdata;
        int_sop      = f0_i1_sop;
        int_eop      = f0_i1_eop;
      end
    default:
      begin
        int_flitdata = {36{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f0_i0_t4_ready = int_ready && (owner == 1'd0);
assign f0_i1_t4_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:36
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:36
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f1_i0
  input  wire            f1_i0_sop,
  input  wire            f1_i0_eop,
  input  wire      [3:0] f1_i0_qos_nxt,
  input  wire      [3:0] f1_i0_qos,
  input  wire     [59:0] f1_i0_flitdata,
  input  wire            f1_i0_t4_activity,
  input  wire            f1_i0_t4_req_nxt,
  input  wire            f1_i0_t4_req,
  output logic           f1_i0_t4_ready,
  // f1_i1
  input  wire            f1_i1_sop,
  input  wire            f1_i1_eop,
  input  wire      [3:0] f1_i1_qos_nxt,
  input  wire      [3:0] f1_i1_qos,
  input  wire     [59:0] f1_i1_flitdata,
  input  wire            f1_i1_t4_activity,
  input  wire            f1_i1_t4_req_nxt,
  input  wire            f1_i1_t4_req,
  output logic           f1_i1_t4_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [59:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [59:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f1_i0_t4_activity || f1_i0_t4_req || f1_i1_t4_activity || f1_i1_t4_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f1_i0_t4_req;
assign nextreqs[0] = f1_i0_t4_req_nxt;
assign nextqos[0] = f1_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f1_i1_t4_req;
assign nextreqs[1] = f1_i1_t4_req_nxt;
assign nextqos[1] = f1_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f1_i0_flitdata;
        int_sop      = f1_i0_sop;
        int_eop      = f1_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f1_i1_flitdata;
        int_sop      = f1_i1_sop;
        int_eop      = f1_i1_eop;
      end
    default:
      begin
        int_flitdata = {60{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f1_i0_t4_ready = int_ready && (owner == 1'd0);
assign f1_i1_t4_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:60
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:60
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_f1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [33:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r0_t4
  output logic           r0_t4_sop,
  output logic           r0_t4_eop,
  output logic     [3:0] r0_t4_qos_nxt,
  output logic     [3:0] r0_t4_qos,
  output logic    [33:0] r0_t4_flitdata,
  output logic           r0_t4_i0_activity,
  output logic           r0_t4_i0_req_nxt,
  output logic           r0_t4_i0_req,
  input  wire            r0_t4_i0_ready,
  output logic           r0_t4_i1_activity,
  output logic           r0_t4_i1_req_nxt,
  output logic           r0_t4_i1_req,
  input  wire            r0_t4_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [33:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [33:0] intp_flitdata;
logic    [33:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:34
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:34
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r0_t4_i0_req = tgtReq[1];
assign tgtXfer[1] = r0_t4_i0_req && r0_t4_i0_ready;
assign r0_t4_i0_activity = tgtAct[1];
assign r0_t4_i0_req_nxt = tgtReqNxt[1];
assign r0_t4_i1_req = tgtReq[0];
assign tgtXfer[0] = r0_t4_i1_req && r0_t4_i1_ready;
assign r0_t4_i1_activity = tgtAct[0];
assign r0_t4_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:34
  .intp_flitdata(intp_flitdata),                                                // o:34
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:34
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r0_t4_sop = intp_sop;
assign r0_t4_eop = intp_eop;
assign r0_t4_qos = intp_qos;
assign r0_t4_flitdata = intp_flitdata;
assign r0_t4_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [33:0] int_flitdata,
  output logic    [33:0] intp_flitdata,
  output logic    [33:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [40:0] wdata;
logic    [40:0] rdata;
logic    [40:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [40:0] fifodata [1:0];
logic    [40:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[35:2] = int_flitdata;
assign intp_flitdata = rdata[35:2];
assign intp_flitdata_nxt = rdata_nxt[35:2];
assign wdata[39:36] = int_qos;
assign intp_qos = rdata[39:36];
assign intp_qos_nxt = rdata_nxt[39:36];
assign wdata[40:40] = int_dstIdx;
assign intp_dstIdx = rdata[40:40];
assign intp_dstIdx_nxt = rdata_nxt[40:40];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {41{1'b0}};
      fifodata[1] <= #1ps {41{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {41{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [23:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r1_t4
  output logic           r1_t4_sop,
  output logic           r1_t4_eop,
  output logic     [3:0] r1_t4_qos_nxt,
  output logic     [3:0] r1_t4_qos,
  output logic    [23:0] r1_t4_flitdata,
  output logic           r1_t4_i0_activity,
  output logic           r1_t4_i0_req_nxt,
  output logic           r1_t4_i0_req,
  input  wire            r1_t4_i0_ready,
  output logic           r1_t4_i1_activity,
  output logic           r1_t4_i1_req_nxt,
  output logic           r1_t4_i1_req,
  input  wire            r1_t4_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [23:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [23:0] intp_flitdata;
logic    [23:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:24
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:24
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r1_t4_i0_req = tgtReq[1];
assign tgtXfer[1] = r1_t4_i0_req && r1_t4_i0_ready;
assign r1_t4_i0_activity = tgtAct[1];
assign r1_t4_i0_req_nxt = tgtReqNxt[1];
assign r1_t4_i1_req = tgtReq[0];
assign tgtXfer[0] = r1_t4_i1_req && r1_t4_i1_ready;
assign r1_t4_i1_activity = tgtAct[0];
assign r1_t4_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:24
  .intp_flitdata(intp_flitdata),                                                // o:24
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:24
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r1_t4_sop = intp_sop;
assign r1_t4_eop = intp_eop;
assign r1_t4_qos = intp_qos;
assign r1_t4_flitdata = intp_flitdata;
assign r1_t4_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [23:0] int_flitdata,
  output logic    [23:0] intp_flitdata,
  output logic    [23:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [30:0] wdata;
logic    [30:0] rdata;
logic    [30:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [30:0] fifodata [1:0];
logic    [30:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[25:2] = int_flitdata;
assign intp_flitdata = rdata[25:2];
assign intp_flitdata_nxt = rdata_nxt[25:2];
assign wdata[29:26] = int_qos;
assign intp_qos = rdata[29:26];
assign intp_qos_nxt = rdata_nxt[29:26];
assign wdata[30:30] = int_dstIdx;
assign intp_dstIdx = rdata[30:30];
assign intp_dstIdx_nxt = rdata_nxt[30:30];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps 31'd0;
      fifodata[1] <= #1ps 31'd0;
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {31{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_usb4_phy_TEA_r1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f0_i0
  input  wire            f0_i0_sop,
  input  wire            f0_i0_eop,
  input  wire      [3:0] f0_i0_qos_nxt,
  input  wire      [3:0] f0_i0_qos,
  input  wire     [35:0] f0_i0_flitdata,
  input  wire            f0_i0_t5_activity,
  input  wire            f0_i0_t5_req_nxt,
  input  wire            f0_i0_t5_req,
  output logic           f0_i0_t5_ready,
  // f0_i1
  input  wire            f0_i1_sop,
  input  wire            f0_i1_eop,
  input  wire      [3:0] f0_i1_qos_nxt,
  input  wire      [3:0] f0_i1_qos,
  input  wire     [35:0] f0_i1_flitdata,
  input  wire            f0_i1_t5_activity,
  input  wire            f0_i1_t5_req_nxt,
  input  wire            f0_i1_t5_req,
  output logic           f0_i1_t5_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [35:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [35:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f0_i0_t5_activity || f0_i0_t5_req || f0_i1_t5_activity || f0_i1_t5_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f0_i0_t5_req;
assign nextreqs[0] = f0_i0_t5_req_nxt;
assign nextqos[0] = f0_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f0_i1_t5_req;
assign nextreqs[1] = f0_i1_t5_req_nxt;
assign nextqos[1] = f0_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f0_i0_flitdata;
        int_sop      = f0_i0_sop;
        int_eop      = f0_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f0_i1_flitdata;
        int_sop      = f0_i1_sop;
        int_eop      = f0_i1_eop;
      end
    default:
      begin
        int_flitdata = {36{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f0_i0_t5_ready = int_ready && (owner == 1'd0);
assign f0_i1_t5_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:36
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:36
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb (
  input  wire            clk,
  input  wire            rst_n,
  // f1_i0
  input  wire            f1_i0_sop,
  input  wire            f1_i0_eop,
  input  wire      [3:0] f1_i0_qos_nxt,
  input  wire      [3:0] f1_i0_qos,
  input  wire     [59:0] f1_i0_flitdata,
  input  wire            f1_i0_t5_activity,
  input  wire            f1_i0_t5_req_nxt,
  input  wire            f1_i0_t5_req,
  output logic           f1_i0_t5_ready,
  // f1_i1
  input  wire            f1_i1_sop,
  input  wire            f1_i1_eop,
  input  wire      [3:0] f1_i1_qos_nxt,
  input  wire      [3:0] f1_i1_qos,
  input  wire     [59:0] f1_i1_flitdata,
  input  wire            f1_i1_t5_activity,
  input  wire            f1_i1_t5_req_nxt,
  input  wire            f1_i1_t5_req,
  output logic           f1_i1_t5_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [59:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [59:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f1_i0_t5_activity || f1_i0_t5_req || f1_i1_t5_activity || f1_i1_t5_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f1_i0_t5_req;
assign nextreqs[0] = f1_i0_t5_req_nxt;
assign nextqos[0] = f1_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f1_i1_t5_req;
assign nextreqs[1] = f1_i1_t5_req_nxt;
assign nextqos[1] = f1_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f1_i0_flitdata;
        int_sop      = f1_i0_sop;
        int_eop      = f1_i0_eop;
      end
    1'd1:
      begin
        int_flitdata = f1_i1_flitdata;
        int_sop      = f1_i1_sop;
        int_eop      = f1_i1_eop;
      end
    default:
      begin
        int_flitdata = {60{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
      end
  endcase
end

// Assign ready bits
assign f1_i0_t5_ready = int_ready && (owner == 1'd0);
assign f1_i1_t5_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:60
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:60
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_f1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [33:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r0_t5
  output logic           r0_t5_sop,
  output logic           r0_t5_eop,
  output logic     [3:0] r0_t5_qos_nxt,
  output logic     [3:0] r0_t5_qos,
  output logic    [33:0] r0_t5_flitdata,
  output logic           r0_t5_i0_activity,
  output logic           r0_t5_i0_req_nxt,
  output logic           r0_t5_i0_req,
  input  wire            r0_t5_i0_ready,
  output logic           r0_t5_i1_activity,
  output logic           r0_t5_i1_req_nxt,
  output logic           r0_t5_i1_req,
  input  wire            r0_t5_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [33:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [33:0] intp_flitdata;
logic    [33:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:34
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:34
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r0_t5_i0_req = tgtReq[1];
assign tgtXfer[1] = r0_t5_i0_req && r0_t5_i0_ready;
assign r0_t5_i0_activity = tgtAct[1];
assign r0_t5_i0_req_nxt = tgtReqNxt[1];
assign r0_t5_i1_req = tgtReq[0];
assign tgtXfer[0] = r0_t5_i1_req && r0_t5_i1_ready;
assign r0_t5_i1_activity = tgtAct[0];
assign r0_t5_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:34
  .intp_flitdata(intp_flitdata),                                                // o:34
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:34
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r0_t5_sop = intp_sop;
assign r0_t5_eop = intp_eop;
assign r0_t5_qos = intp_qos;
assign r0_t5_flitdata = intp_flitdata;
assign r0_t5_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [33:0] int_flitdata,
  output logic    [33:0] intp_flitdata,
  output logic    [33:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [40:0] wdata;
logic    [40:0] rdata;
logic    [40:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [40:0] fifodata [1:0];
logic    [40:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[35:2] = int_flitdata;
assign intp_flitdata = rdata[35:2];
assign intp_flitdata_nxt = rdata_nxt[35:2];
assign wdata[39:36] = int_qos;
assign intp_qos = rdata[39:36];
assign intp_qos_nxt = rdata_nxt[39:36];
assign wdata[40:40] = int_dstIdx;
assign intp_dstIdx = rdata[40:40];
assign intp_dstIdx_nxt = rdata_nxt[40:40];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {41{1'b0}};
      fifodata[1] <= #1ps {41{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {41{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec (
  input  wire            clk,
  input  wire            rst_n,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [23:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r1_t5
  output logic           r1_t5_sop,
  output logic           r1_t5_eop,
  output logic     [3:0] r1_t5_qos_nxt,
  output logic     [3:0] r1_t5_qos,
  output logic    [23:0] r1_t5_flitdata,
  output logic           r1_t5_i0_activity,
  output logic           r1_t5_i0_req_nxt,
  output logic           r1_t5_i0_req,
  input  wire            r1_t5_i0_ready,
  output logic           r1_t5_i1_activity,
  output logic           r1_t5_i1_req_nxt,
  output logic           r1_t5_i1_req,
  input  wire            r1_t5_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [23:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [23:0] intp_flitdata;
logic    [23:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [2:0] int_destid;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic     [0:0] tmp_dstIdx;
logic     [0:0] int_dstIdx;
logic     [0:0] dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:24
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:24
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? dstIdx : intp_dstIdx;
assign int_destid = int_flitdata[3+3:4];
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r1_t5_i0_req = tgtReq[1];
assign tgtXfer[1] = r1_t5_i0_req && r1_t5_i0_ready;
assign r1_t5_i0_activity = tgtAct[1];
assign r1_t5_i0_req_nxt = tgtReqNxt[1];
assign r1_t5_i1_req = tgtReq[0];
assign tgtXfer[0] = r1_t5_i1_req && r1_t5_i1_ready;
assign r1_t5_i1_activity = tgtAct[0];
assign r1_t5_i1_req_nxt = tgtReqNxt[0];
assign tmp_dstIdx[0] = ((int_destid == 3'd1));
assign int_dstIdx = tmp_dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:24
  .intp_flitdata(intp_flitdata),                                                // o:24
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:24
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r1_t5_sop = intp_sop;
assign r1_t5_eop = intp_eop;
assign r1_t5_qos = intp_qos;
assign r1_t5_flitdata = intp_flitdata;
assign r1_t5_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [23:0] int_flitdata,
  output logic    [23:0] intp_flitdata,
  output logic    [23:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [30:0] wdata;
logic    [30:0] rdata;
logic    [30:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [30:0] fifodata [1:0];
logic    [30:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[25:2] = int_flitdata;
assign intp_flitdata = rdata[25:2];
assign intp_flitdata_nxt = rdata_nxt[25:2];
assign wdata[29:26] = int_qos;
assign intp_qos = rdata[29:26];
assign intp_qos_nxt = rdata_nxt[29:26];
assign wdata[30:30] = int_dstIdx;
assign intp_dstIdx = rdata[30:30];
assign intp_dstIdx_nxt = rdata_nxt[30:30];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps 31'd0;
      fifodata[1] <= #1ps 31'd0;
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {31{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_pam3_xcvr_TEA_r1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f0_arb (
  input  wire            clk,
  input  wire            rst_n,
  output logic     [0:0] srcIdx,
  // f0_i0
  input  wire            f0_i0_sop,
  input  wire            f0_i0_eop,
  input  wire      [3:0] f0_i0_qos_nxt,
  input  wire      [3:0] f0_i0_qos,
  input  wire     [35:0] f0_i0_flitdata,
  input  wire            f0_i0_t1000_activity,
  input  wire            f0_i0_t1000_req_nxt,
  input  wire            f0_i0_t1000_req,
  output logic           f0_i0_t1000_ready,
  // f0_i1
  input  wire            f0_i1_sop,
  input  wire            f0_i1_eop,
  input  wire      [3:0] f0_i1_qos_nxt,
  input  wire      [3:0] f0_i1_qos,
  input  wire     [35:0] f0_i1_flitdata,
  input  wire            f0_i1_t1000_activity,
  input  wire            f0_i1_t1000_req_nxt,
  input  wire            f0_i1_t1000_req,
  output logic           f0_i1_t1000_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [35:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [35:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f0_i0_t1000_activity || f0_i0_t1000_req || f0_i1_t1000_activity || f0_i1_t1000_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_t1000_f0_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f0_i0_t1000_req;
assign nextreqs[0] = f0_i0_t1000_req_nxt;
assign nextqos[0] = f0_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f0_i1_t1000_req;
assign nextreqs[1] = f0_i1_t1000_req_nxt;
assign nextqos[1] = f0_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f0_i0_flitdata;
        int_sop      = f0_i0_sop;
        int_eop      = f0_i0_eop;
        srcIdx       = 1'd0;
      end
    1'd1:
      begin
        int_flitdata = f0_i1_flitdata;
        int_sop      = f0_i1_sop;
        int_eop      = f0_i1_eop;
        srcIdx       = 1'd1;
      end
    default:
      begin
        int_flitdata = {36{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
        srcIdx       = 1'd0;
      end
  endcase
end

// Assign ready bits
assign f0_i0_t1000_ready = int_ready && (owner == 1'd0);
assign f0_i1_t1000_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_t1000_f0_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:36
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:36
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f0_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f0_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_t1000_f0_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f0_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f1_arb (
  input  wire            clk,
  input  wire            rst_n,
  output logic     [0:0] srcIdx,
  // f1_i0
  input  wire            f1_i0_sop,
  input  wire            f1_i0_eop,
  input  wire      [3:0] f1_i0_qos_nxt,
  input  wire      [3:0] f1_i0_qos,
  input  wire     [59:0] f1_i0_flitdata,
  input  wire            f1_i0_t1000_activity,
  input  wire            f1_i0_t1000_req_nxt,
  input  wire            f1_i0_t1000_req,
  output logic           f1_i0_t1000_ready,
  // f1_i1
  input  wire            f1_i1_sop,
  input  wire            f1_i1_eop,
  input  wire      [3:0] f1_i1_qos_nxt,
  input  wire      [3:0] f1_i1_qos,
  input  wire     [59:0] f1_i1_flitdata,
  input  wire            f1_i1_t1000_activity,
  input  wire            f1_i1_t1000_req_nxt,
  input  wire            f1_i1_t1000_req,
  output logic           f1_i1_t1000_ready,
  // tgt
  output logic           tgt_activity,                                          // Upcoming activity indicator
  output logic           tgt_req,                                               // Flit transfer request
  output logic           tgt_sop,                                               // Start of packet indicator
  output logic           tgt_eop,                                               // End of packet indicator
  output logic    [59:0] tgt_flitdata,                                          // Flit data
  input  wire            tgt_ready                                              // Flit transfer ready
);

logic           int_activity;
logic           int_req;
logic           int_ready;
logic    [59:0] int_flitdata;
logic           int_sop;
logic           int_eop;
logic     [0:0] int_vc;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [0:0] owner;                                                          // This is the new owner when arbitration occurrs
logic           rearbitrate;                                                    // This signal indicates that arbitration is happening
logic     [1:0] prawreqs;                                                       // Raw reqs are the req signals from the decoder
logic     [1:0] nextreqs;                                                       // Next reqs are the req signals coming up next cycle
logic     [1:0] preqs;                                                          // preqs are verified arbitration candidates
logic     [4:0] nextqos [1:0];                                                  // Next QOS are next qos values scaled by 1 to be 1 to 16.
logic     [4:0] tscore [1:0];
logic     [4:0] tscore_nxt [1:0];
logic     [1:0] tscore_en;
logic     [0:0] powner;
logic     [4:0] maxScore;
logic     [4:0] maxScore_nxt;
logic     [0:0] maxScore_en;
logic     [4:0] tmpMax0;
logic     [0:0] busy;
logic     [0:0] busy_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Interface to Decoders
// ============================================================================
// ============================================================================
// Target Port Interface
// ============================================================================
assign frst_n = rst_n;
assign int_activity = f1_i0_t1000_activity || f1_i0_t1000_req || f1_i1_t1000_activity || f1_i1_t1000_req;
// Data Array Clock Gating Logic
assign gclkEn = int_activity;
usb4_tc_noc_rtr0_t1000_f1_arb_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// tscore is the total score of the channel, capped to 0x1F
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      tscore[0] <= #1ps 5'd0;
      tscore[1] <= #1ps 5'd0;
    end
  else
    begin
      if (tscore_en[0])
        tscore[0] <= #1ps tscore_nxt[0];
      if (tscore_en[1])
        tscore[1] <= #1ps tscore_nxt[1];
    end
end

// powner is the last successful arbitrated channel number
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    powner <= #1ps 1'd0;
  else if (int_req)
    powner <= #1ps owner;
end

// maxScore is the highest score of all channels
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    maxScore <= #1ps 5'd0;
  else if (maxScore_en)
    maxScore <= #1ps maxScore_nxt;
end

assign prawreqs[0] = f1_i0_t1000_req;
assign nextreqs[0] = f1_i0_t1000_req_nxt;
assign nextqos[0] = f1_i0_qos_nxt + 4'd1;
assign prawreqs[1] = f1_i1_t1000_req;
assign nextreqs[1] = f1_i1_t1000_req_nxt;
assign nextqos[1] = f1_i1_qos_nxt + 4'd1;
// Bump tscore for next cycle.
always_comb
begin
    tscore_nxt[0] = tscore[0];
    tscore_nxt[1] = tscore[1];
    tscore_en  = 2'd0;
    if( rearbitrate )
      begin
        // Processing in an Arbitration Cycle
        // If this channel was selected or is idle, score it zero
        // Else if score == 0, then start off with rawqos
        // Else if not capped at 0x1F, bump it
        tscore_en  = {2{1'b1}};
        if( owner==1'd0 || tscore[0] == 5'd0 )
          tscore_nxt[0] = nextreqs[0] ? nextqos[0] : 5'd0;
        else if( tscore[0]!=5'h1F )
          tscore_nxt[0] = tscore[0]+5'd1;
        if( owner==1'd1 || tscore[1] == 5'd0 )
          tscore_nxt[1] = nextreqs[1] ? nextqos[1] : 5'd0;
        else if( tscore[1]!=5'h1F )
          tscore_nxt[1] = tscore[1]+5'd1;
      end
    else
      begin
        // Processing for a non-Arbitration Cycle
        // If score is zero and channel is requesting, start off with rawqos
        if( tscore[0] == 5'd0 && nextreqs[0] && (!busy || powner != 1'd0) )
          begin
            tscore_en[0]  = 1'b1;
            tscore_nxt[0] = nextqos[0];
          end
        if( tscore[1] == 5'd0 && nextreqs[1] && (!busy || powner != 1'd1) )
          begin
            tscore_en[1]  = 1'b1;
            tscore_nxt[1] = nextqos[1];
          end
      end
end

// Code to find the highest score of any requestor
assign tmpMax0 = tscore_nxt[1]>tscore_nxt[0] ? tscore_nxt[1] : tscore_nxt[0];
assign maxScore_nxt = tmpMax0;
assign maxScore_en = 1'b1;
// Any request from a channel at maxScore is filtered through
always_comb
begin
  preqs = 2'd0;
  if( tscore[0]==maxScore )
    preqs[0] = prawreqs[0];
  if( tscore[1]==maxScore )
    preqs[1] = prawreqs[1];
end

// Find highest priority requester in priority tier $pri based on previous owner
always_comb
begin
  if (busy)
    begin
      owner = powner;
    end
  else
    begin
      case (powner)
        1'd0: owner = (preqs[1]) ? 1'd1 :  powner;
        1'd1: owner = (preqs[0]) ? 1'd0 :  powner;
        default: owner = powner;
      endcase
    end
end

// Target request is asserted anytime any initiator is requesting when not busy
// but only when specific request corresponding to current owner when busy
assign int_req = (busy) ? prawreqs[owner] : |preqs;
// Signal which indicates its time to rearbitrate
assign rearbitrate = int_req && !busy_nxt;
// Mux output signals
always_comb
begin
  case(owner)
    1'd0:
      begin
        int_flitdata = f1_i0_flitdata;
        int_sop      = f1_i0_sop;
        int_eop      = f1_i0_eop;
        srcIdx       = 1'd0;
      end
    1'd1:
      begin
        int_flitdata = f1_i1_flitdata;
        int_sop      = f1_i1_sop;
        int_eop      = f1_i1_eop;
        srcIdx       = 1'd1;
      end
    default:
      begin
        int_flitdata = {60{1'b0}};
        int_sop      = 1'b0;
        int_eop      = 1'b0;
        srcIdx       = 1'd0;
      end
  endcase
end

// Assign ready bits
assign f1_i0_t1000_ready = int_ready && (owner == 1'd0);
assign f1_i1_t1000_ready = int_ready && (owner == 1'd1);
// Arbiter busy indicator
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    busy <= #1ps 1'd0;
  else
    busy <= #1ps busy_nxt;
end

always_comb
begin
  busy_nxt = busy;
  if (int_req && int_ready && int_eop)
    busy_nxt = 1'b0;
  else if (int_req)
    busy_nxt = 1'b1;
end

// ============================================================================
// Target Port $i Egress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_t1000_f1_arb_ep ep (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(int_activity),                                                  // i:1
  .src_req(int_req),                                                            // i:1
  .src_sop(int_sop),                                                            // i:1
  .src_eop(int_eop),                                                            // i:1
  .src_flitdata(int_flitdata),                                                  // i:60
  .src_ready(int_ready),                                                        // o:1
  .dst_activity(tgt_activity),                                                  // o:1
  .dst_req(tgt_req),                                                            // o:1
  .dst_sop(tgt_sop),                                                            // o:1
  .dst_eop(tgt_eop),                                                            // o:1
  .dst_flitdata(tgt_flitdata),                                                  // o:60
  .dst_ready(tgt_ready)                                                         // i:1
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f1_arb_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f1_arb_ep (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_t1000_f1_arb_ep_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_f1_arb_ep_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r0_dec (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [0:0] dstIdx,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [33:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r0_t1000
  output logic           r0_t1000_sop,
  output logic           r0_t1000_eop,
  output logic     [3:0] r0_t1000_qos_nxt,
  output logic     [3:0] r0_t1000_qos,
  output logic    [33:0] r0_t1000_flitdata,
  output logic           r0_t1000_i0_activity,
  output logic           r0_t1000_i0_req_nxt,
  output logic           r0_t1000_i0_req,
  input  wire            r0_t1000_i0_ready,
  output logic           r0_t1000_i1_activity,
  output logic           r0_t1000_i1_req_nxt,
  output logic           r0_t1000_i1_req,
  input  wire            r0_t1000_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [33:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [33:0] intp_flitdata;
logic    [33:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic           int_inPkt;
logic     [0:0] int_dstIdx;
logic     [0:0] held_dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_t1000_r0_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:34
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:34
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_t1000_r0_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

assign int_inPkt = inPkt;
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    held_dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    held_dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? held_dstIdx : intp_dstIdx;
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r0_t1000_i0_req = tgtReq[0];
assign tgtXfer[0] = r0_t1000_i0_req && r0_t1000_i0_ready;
assign r0_t1000_i0_activity = tgtAct[0];
assign r0_t1000_i0_req_nxt = tgtReqNxt[0];
assign r0_t1000_i1_req = tgtReq[1];
assign tgtXfer[1] = r0_t1000_i1_req && r0_t1000_i1_ready;
assign r0_t1000_i1_activity = tgtAct[1];
assign r0_t1000_i1_req_nxt = tgtReqNxt[1];
assign int_dstIdx = dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_t1000_r0_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:34
  .intp_flitdata(intp_flitdata),                                                // o:34
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:34
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r0_t1000_sop = intp_sop;
assign r0_t1000_eop = intp_eop;
assign r0_t1000_qos = intp_qos;
assign r0_t1000_flitdata = intp_flitdata;
assign r0_t1000_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r0_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_t1000_r0_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r0_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r0_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r0_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [33:0] int_flitdata,
  output logic    [33:0] intp_flitdata,
  output logic    [33:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [40:0] wdata;
logic    [40:0] rdata;
logic    [40:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [40:0] fifodata [1:0];
logic    [40:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_t1000_r0_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[35:2] = int_flitdata;
assign intp_flitdata = rdata[35:2];
assign intp_flitdata_nxt = rdata_nxt[35:2];
assign wdata[39:36] = int_qos;
assign intp_qos = rdata[39:36];
assign intp_qos_nxt = rdata_nxt[39:36];
assign wdata[40:40] = int_dstIdx;
assign intp_dstIdx = rdata[40:40];
assign intp_dstIdx_nxt = rdata_nxt[40:40];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps {41{1'b0}};
      fifodata[1] <= #1ps {41{1'b0}};
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {41{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r0_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r1_dec (
  input  wire            clk,
  input  wire            rst_n,
  input  wire      [0:0] dstIdx,
  // ini
  input  wire            ini_activity,                                          // Upcoming activity indicator
  input  wire            ini_req,                                               // Flit transfer request
  input  wire            ini_sop,                                               // Start of packet indicator
  input  wire            ini_eop,                                               // End of packet indicator
  input  wire     [23:0] ini_flitdata,                                          // Flit data
  output logic           ini_ready,                                             // Flit transfer ready
  // r1_t1000
  output logic           r1_t1000_sop,
  output logic           r1_t1000_eop,
  output logic     [3:0] r1_t1000_qos_nxt,
  output logic     [3:0] r1_t1000_qos,
  output logic    [23:0] r1_t1000_flitdata,
  output logic           r1_t1000_i0_activity,
  output logic           r1_t1000_i0_req_nxt,
  output logic           r1_t1000_i0_req,
  input  wire            r1_t1000_i0_ready,
  output logic           r1_t1000_i1_activity,
  output logic           r1_t1000_i1_req_nxt,
  output logic           r1_t1000_i1_req,
  input  wire            r1_t1000_i1_ready
);

logic           int_activity;                                                   // Upcoming activity indicator
logic           int_req;                                                        // Flit transfer request
logic           int_sop;                                                        // Start of packet indicator
logic           int_eop;                                                        // End of packet indicator
logic    [23:0] int_flitdata;                                                   // Flit data
logic           int_ready;                                                      // Flit transfer ready
logic           intp_sop;
logic           intp_sop_nxt;
logic           intp_eop;
logic           intp_eop_nxt;
logic    [23:0] intp_flitdata;
logic    [23:0] intp_flitdata_nxt;
logic     [3:0] intp_qos;
logic     [3:0] intp_qos_nxt;
logic           intp_dstIdx;
logic           intp_dstIdx_nxt;
logic           frst_n;
logic           gclk;
wire            gclkEn;
wire            gclkAct;
logic     [3:0] qos;
logic     [3:0] int_qos;
logic     [0:0] inPkt;
logic           int_inPkt;
logic     [0:0] int_dstIdx;
logic     [0:0] held_dstIdx;
logic     [0:0] useDstIdx;
logic     [1:0] tgtReq;
logic     [1:0] tgtAct;
logic     [1:0] tgtXfer;
logic     [1:0] tgtReqNxt;
logic     [1:0] lockedDest;
logic           intp_ready;
logic           intp_req;
logic           intp_activity;
logic           intp_req_nxt;
// ============================================================================
// Clock and reset
// ============================================================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================================================
// Initiator  Interface (LLK subordinate)
// ============================================================================
// ============================================================================
// Interface to Arbiters
// ============================================================================
// ============================================================================
// Ingress Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_t1000_r1_dec_ip ip (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ini_activity),                                                  // i:1
  .src_req(ini_req),                                                            // i:1
  .src_sop(ini_sop),                                                            // i:1
  .src_eop(ini_eop),                                                            // i:1
  .src_flitdata(ini_flitdata),                                                  // i:24
  .src_ready(ini_ready),                                                        // o:1
  .dst_activity(int_activity),                                                  // o:1
  .dst_req(int_req),                                                            // o:1
  .dst_sop(int_sop),                                                            // o:1
  .dst_eop(int_eop),                                                            // o:1
  .dst_flitdata(int_flitdata),                                                  // o:24
  .dst_ready(int_ready)                                                         // i:1
);
assign frst_n = rst_n;
// ============================================================================
// Clock Gating
// ============================================================================
// Data Array Clock Gating Logic
assign gclkEn = int_activity || intp_activity || int_req || intp_req;
usb4_tc_noc_rtr0_t1000_r1_dec_cg cg (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .enbIn(gclkEn),                                                               // i:1
  .clkOut(gclk),                                                                // o:1
  .isActive(gclkAct)                                                            // o:1
);
// Pipe Ingress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    qos <= #1ps 4'd0;
  else if (int_req && int_ready && int_sop)
    qos <= #1ps int_flitdata[3:0];
end

assign int_qos = int_sop ? int_flitdata[3:0] : qos;
// Pipe Egress Flops
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    inPkt <= #1ps 1'd0;
  else if (intp_req && intp_ready)
    inPkt <= #1ps ~intp_eop;
end

assign int_inPkt = inPkt;
always_ff @(posedge gclk, negedge frst_n)
begin
  if (!frst_n)
    held_dstIdx <= #1ps 1'd0;
  else if (intp_req && intp_ready && intp_sop)
    held_dstIdx <= #1ps intp_dstIdx;
end

assign useDstIdx = inPkt ? held_dstIdx : intp_dstIdx;
// ============================================================================
// Perform the actual decode of the destination ID
// ============================================================================
assign r1_t1000_i0_req = tgtReq[0];
assign tgtXfer[0] = r1_t1000_i0_req && r1_t1000_i0_ready;
assign r1_t1000_i0_activity = tgtAct[0];
assign r1_t1000_i0_req_nxt = tgtReqNxt[0];
assign r1_t1000_i1_req = tgtReq[1];
assign tgtXfer[1] = r1_t1000_i1_req && r1_t1000_i1_ready;
assign r1_t1000_i1_activity = tgtAct[1];
assign r1_t1000_i1_req_nxt = tgtReqNxt[1];
assign int_dstIdx = dstIdx;
assign lockedDest = 2'd1 << useDstIdx;
always_comb
begin
  tgtReq = 2'd0;
  if( intp_req )
    tgtReq = lockedDest;
end

always_comb
begin
  tgtAct = 2'd0;
  if( intp_activity || (int_activity && !inPkt) )
    begin
      if( !inPkt || (intp_req && intp_eop) )
        tgtAct = {2{1'b1}};
      else
        tgtAct = lockedDest;
    end
end

always_comb
begin
  tgtReqNxt = 2'd0;
  if( intp_req_nxt )
    begin
      if( intp_sop_nxt )
        tgtReqNxt = 2'd1 << intp_dstIdx_nxt;
      else
        tgtReqNxt = lockedDest;
    end
end

// ============================================================================
// Center Pipe Stage
// ============================================================================
usb4_tc_noc_rtr0_t1000_r1_dec_cp cp (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(int_req),                                                               // i:1
  .wact(int_activity),                                                          // i:1
  .ract(intp_activity),                                                         // o:1
  .wrdy(int_ready),                                                             // o:1
  .rreq(intp_ready),                                                            // i:1
  .rrdy(intp_req),                                                              // o:1
  .rrdy_nxt(intp_req_nxt),                                                      // o:1
  .int_sop(int_sop),                                                            // i:1
  .intp_sop(intp_sop),                                                          // o:1
  .intp_sop_nxt(intp_sop_nxt),                                                  // o:1
  .int_eop(int_eop),                                                            // i:1
  .intp_eop(intp_eop),                                                          // o:1
  .intp_eop_nxt(intp_eop_nxt),                                                  // o:1
  .int_flitdata(int_flitdata),                                                  // i:24
  .intp_flitdata(intp_flitdata),                                                // o:24
  .intp_flitdata_nxt(intp_flitdata_nxt),                                        // o:24
  .int_qos(int_qos),                                                            // i:4
  .intp_qos(intp_qos),                                                          // o:4
  .intp_qos_nxt(intp_qos_nxt),                                                  // o:4
  .int_dstIdx(int_dstIdx),                                                      // i:1
  .intp_dstIdx(intp_dstIdx),                                                    // o:1
  .intp_dstIdx_nxt(intp_dstIdx_nxt)                                             // o:1
);
// Pop the center pipeline stage
assign intp_ready = tgtXfer[useDstIdx];
// Assign the remaining outputs
assign r1_t1000_sop = intp_sop;
assign r1_t1000_eop = intp_eop;
assign r1_t1000_qos = intp_qos;
assign r1_t1000_flitdata = intp_flitdata;
assign r1_t1000_qos_nxt = intp_qos_nxt;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r1_dec_ip (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_t1000_r1_dec_ip_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r1_dec_ip_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r1_dec_cg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r1_dec_cp (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  output logic           rrdy_nxt,
  input  wire            int_sop,
  output logic           intp_sop,
  output logic           intp_sop_nxt,
  input  wire            int_eop,
  output logic           intp_eop,
  output logic           intp_eop_nxt,
  input  wire     [23:0] int_flitdata,
  output logic    [23:0] intp_flitdata,
  output logic    [23:0] intp_flitdata_nxt,
  input  wire      [3:0] int_qos,
  output logic     [3:0] intp_qos,
  output logic     [3:0] intp_qos_nxt,
  input  wire            int_dstIdx,
  output logic           intp_dstIdx,
  output logic           intp_dstIdx_nxt
);

logic           valid_wr;
logic           valid_rd;
logic    [30:0] wdata;
logic    [30:0] rdata;
logic    [30:0] rdata_nxt;
logic           cclk;
logic           dclk;
logic           dclkAct;
logic           cclkAct;
wire            dclkEn;
logic     [0:0] d1wact;
logic     [0:0] wptr;
logic     [0:0] wptr_nxt;
logic     [0:0] wptr_en;
logic    [30:0] fifodata [1:0];
logic    [30:0] fifodata_nxt [1:0];
logic     [1:0] fifodata_en;
logic     [0:0] rptr;
logic     [0:0] rptr_nxt;
logic     [0:0] rptr_en;
logic     [1:0] occ;
logic     [1:0] occ_nxt;
logic     [0:0] occ_en;
logic     [0:0] iwrdy;
logic     [0:0] iwrdy_nxt;
logic     [0:0] iwrdy_en;
logic     [0:0] irrdy;
logic     [0:0] irrdy_nxt;
assign valid_wr = wreq && wrdy;
assign valid_rd = rreq && rrdy;
// ==============================================
// Power Management Control
// ==============================================
// Data Array Clock Gating Logic
assign dclkEn = wreq || wact || (|occ);
usb4_tc_noc_rtr0_t1000_r1_dec_cp_dcg dcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(dclkEn),                                                               // i:1
  .clkOut(dclk),                                                                // o:1
  .isActive(dclkAct)                                                            // o:1
);
// Control Signals Clock Gating Logic
assign cclk = dclk;
assign cclkAct = dclkAct;
// wire  cclkEn = wreq || wact || |occ;
// minst clockGate ccg ( #arst($arst) #regEnable(1) #inclTMode($inclTMode) #idleWait(0) .*(*) .clk(clk) .rst_n(rst_n) .enbIn(cclkEn) .clkOut(cclk) .isActive(cclkAct));
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    d1wact <= #1ps 1'd0;
  else
    d1wact <= #1ps wreq || wact;
end

assign ract = d1wact || irrdy || irrdy_nxt;
assign wdata[0:0] = int_sop;
assign intp_sop = rdata[0:0];
assign intp_sop_nxt = rdata_nxt[0:0];
assign wdata[1:1] = int_eop;
assign intp_eop = rdata[1:1];
assign intp_eop_nxt = rdata_nxt[1:1];
assign wdata[25:2] = int_flitdata;
assign intp_flitdata = rdata[25:2];
assign intp_flitdata_nxt = rdata_nxt[25:2];
assign wdata[29:26] = int_qos;
assign intp_qos = rdata[29:26];
assign intp_qos_nxt = rdata_nxt[29:26];
assign wdata[30:30] = int_dstIdx;
assign intp_dstIdx = rdata[30:30];
assign intp_dstIdx_nxt = rdata_nxt[30:30];
// Write pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    wptr <= #1ps 1'd0;
  else if (wptr_en)
    wptr <= #1ps wptr_nxt;
end

always_comb
begin
  wptr_nxt = wptr;
  wptr_en = 1'b0;
  if (valid_wr && (wptr == 1'd1))
    begin
      wptr_nxt = 1'd0;
      wptr_en  = 1'b1;
    end
  else if (valid_wr)
    begin
      wptr_nxt = wptr + 1'd1;
      wptr_en  = 1'b1;
    end
end

// Write data
always_ff @(posedge dclk, negedge rst_n)
begin
  if (!rst_n)
    begin
      fifodata[0] <= #1ps 31'd0;
      fifodata[1] <= #1ps 31'd0;
    end
  else
    begin
      if (fifodata_en[0])
        fifodata[0] <= #1ps fifodata_nxt[0];
      if (fifodata_en[1])
        fifodata[1] <= #1ps fifodata_nxt[1];
    end
end

always_comb
begin
  fifodata_nxt[0] = fifodata[0];
  fifodata_nxt[1] = fifodata[1];
  fifodata_en  = {2{1'b0}};
  if (valid_wr)
    begin
      fifodata_nxt[wptr] = wdata;
      fifodata_en[wptr]  = 1'b1;
    end
end

// Read Pointer
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    rptr <= #1ps 1'd0;
  else if (rptr_en)
    rptr <= #1ps rptr_nxt;
end

always_comb
begin
  rptr_nxt = rptr;
  rptr_en  = 1'b0;
  if (valid_rd && (rptr == 1'd1))
    begin
      rptr_nxt       = 1'd0;
      rptr_en        = 1'b1;
    end
  else if (valid_rd)
    begin
      rptr_nxt       = rptr + 1'd1;
      rptr_en        = 1'b1;
    end
end

// Occupancy
always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    occ <= #1ps 2'd0;
  else if (occ_en)
    occ <= #1ps occ_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    iwrdy <= #1ps 1'b0;
  else if (iwrdy_en)
    iwrdy <= #1ps iwrdy_nxt;
end

always_ff @(posedge cclk, negedge rst_n)
begin
  if (!rst_n)
    irrdy <= #1ps 1'd0;
  else if (occ_en)
    irrdy <= #1ps irrdy_nxt;
end

always_comb
begin
  occ_nxt   = occ;
  iwrdy_nxt = iwrdy;
  irrdy_nxt = irrdy;
  occ_en    = 1'b0;
  iwrdy_en  = 1'b0;
  if (valid_wr && !valid_rd)
    begin
      occ_nxt   = occ + 2'd1;
      iwrdy_nxt = (occ < 2'd1);
      irrdy_nxt = 1'b1;
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!valid_wr && valid_rd)
    begin
      occ_nxt   = occ - 2'd1;
      iwrdy_nxt = 1'b1;
      irrdy_nxt = (occ > 2'd1);
      occ_en    = 1'b1;
      iwrdy_en  = 1'b1;
    end
  else if (!iwrdy && occ < 2'd1)
    begin
      iwrdy_nxt = 1'b1;
      iwrdy_en  = 1'b1;
    end
end

// Create the external ready signals based on internal signals and clock run state
assign wrdy = iwrdy && cclkAct && dclkAct;
assign rrdy = irrdy && cclkAct;
// Read data
assign rdata = fifodata[rptr];
assign rrdy_nxt = irrdy_nxt;
assign rdata_nxt = irrdy_nxt ? fifodata_nxt[rptr_nxt] : {31{1'b0}};
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_t1000_r1_dec_cp_dcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt (
  input  wire            clk,
  input  wire            rst_n,
  output logic           regWReq,
  output logic     [9:0] regWAddr,
  output logic    [31:0] regWData,
  output logic     [3:0] regWEn,
  output logic           regRReq,
  output logic     [9:0] regRAddr,
  input  wire     [31:0] regRData,
  input  wire      [0:0] f0_srcIdx,
  input  wire      [0:0] f1_srcIdx,
  output wire      [0:0] r0_dstIdx,
  output wire      [0:0] r1_dstIdx,
  // f0
  input  wire            f0_activity,                                           // Upcoming activity indicator
  input  wire            f0_req,                                                // Flit transfer request
  input  wire            f0_sop,                                                // Start of packet indicator
  input  wire            f0_eop,                                                // End of packet indicator
  input  wire     [35:0] f0_flitdata,                                           // Flit data
  output logic           f0_ready,                                              // Flit transfer ready
  // f1
  input  wire            f1_activity,                                           // Upcoming activity indicator
  input  wire            f1_req,                                                // Flit transfer request
  input  wire            f1_sop,                                                // Start of packet indicator
  input  wire            f1_eop,                                                // End of packet indicator
  input  wire     [59:0] f1_flitdata,                                           // Flit data
  output logic           f1_ready,                                              // Flit transfer ready
  // r0
  output logic           r0_activity,                                           // Upcoming activity indicator
  output logic           r0_req,                                                // Flit transfer request
  output logic           r0_sop,                                                // Start of packet indicator
  output logic           r0_eop,                                                // End of packet indicator
  output logic    [33:0] r0_flitdata,                                           // Flit data
  input  wire            r0_ready,                                              // Flit transfer ready
  // r1
  output logic           r1_activity,                                           // Upcoming activity indicator
  output logic           r1_req,                                                // Flit transfer request
  output logic           r1_sop,                                                // Start of packet indicator
  output logic           r1_eop,                                                // End of packet indicator
  output logic    [23:0] r1_flitdata,                                           // Flit data
  input  wire            r1_ready                                               // Flit transfer ready
);

logic           if0_activity;                                                   // Upcoming activity indicator
logic           if0_req;                                                        // Flit transfer request
logic           if0_sop;                                                        // Start of packet indicator
logic           if0_eop;                                                        // End of packet indicator
logic    [35:0] if0_flitdata;                                                   // Flit data
logic           if0_ready;                                                      // Flit transfer ready
logic           if1_activity;                                                   // Upcoming activity indicator
logic           if1_req;                                                        // Flit transfer request
logic           if1_sop;                                                        // Start of packet indicator
logic           if1_eop;                                                        // End of packet indicator
logic    [59:0] if1_flitdata;                                                   // Flit data
logic           if1_ready;                                                      // Flit transfer ready
logic           ir0_activity;                                                   // Upcoming activity indicator
logic           ir0_req;                                                        // Flit transfer request
logic           ir0_sop;                                                        // Start of packet indicator
logic           ir0_eop;                                                        // End of packet indicator
logic    [33:0] ir0_flitdata;                                                   // Flit data
logic           ir0_ready;                                                      // Flit transfer ready
logic           ir1_activity;                                                   // Upcoming activity indicator
logic           ir1_req;                                                        // Flit transfer request
logic           ir1_sop;                                                        // Start of packet indicator
logic           ir1_eop;                                                        // End of packet indicator
logic    [23:0] ir1_flitdata;                                                   // Flit data
logic           ir1_ready;                                                      // Flit transfer ready
logic    [23:0] ws_hdr;                                                         // Packed header
logic           wc_buf_we;
logic    [71:0] wc_bus;
logic     [2:0] int_awsid;
logic     [2:0] int_awdid;
logic     [1:0] int_awid;
logic     [3:0] int_awqos;
logic     [1:0] int_awbar;
logic    [67:0] rds_hdr;
logic           rc_buf_we;
logic    [59:0] rc_bus;
logic           frst_n;
logic           wclk;
wire            wclkEn;
logic           rclk;
wire            rclkEn;
logic     [0:0] wc_cnt;
logic     [0:0] wc_cnt_nxt;
logic     [0:0] wc_cnt_en;
logic     [0:0] wr_portIdx;
logic     [0:0] wr_portIdx_nxt;
logic     [0:0] wr_portIdx_en;
logic     [0:0] ws_cnt;
logic     [0:0] ws_cnt_nxt;
logic     [0:0] ws_cnt_en;
logic     [1:0] wcd_state;
logic     [1:0] wcd_state_nxt;
logic     [0:0] wcd_state_en;
logic    [35:0] wc_buf [1:0];
logic     [1:0] wc_buf_en;
logic    [35:0] wregdata;
logic    [35:0] wregdata_nxt;
logic     [0:0] wregdata_en;
logic     [1:0] wregmode;
logic     [1:0] wregmode_nxt;
logic     [0:0] wregmode_en;
logic    [31:0] writeAddr;
logic     [0:0] segIdx;
logic    [35:0] flitSeg [0:0];
logic     [0:0] rc_cnt;
logic     [0:0] rc_cnt_nxt;
logic     [0:0] rc_cnt_en;
logic    [59:0] rc_buf [0:0];
logic     [0:0] rc_buf_en;
logic     [0:0] rc_portIdx;
logic     [0:0] rc_portIdx_nxt;
logic     [0:0] rc_portIdx_en;
logic           int_arIsCMO;
logic     [2:0] int_rplen;
logic    [31:0] int_araddr;
logic     [2:0] int_ardid;
logic           isNarrow;
logic     [0:0] rds_cnt;
logic     [0:0] rds_cnt_nxt;
logic     [0:0] rds_cnt_en;
logic     [1:0] rds_state;
logic     [1:0] rds_state_nxt;
logic     [0:0] rds_state_en;
logic     [8:0] oLoop;
logic     [8:0] oLoop_nxt;
logic     [0:0] oLoop_en;
logic     [5:0] iLoop;
logic     [5:0] iLoop_nxt;
logic     [0:0] iLoop_en;
logic     [3:0] int_arsize;
logic     [1:0] int_arburst;
logic     [3:0] tmp_arsize;
logic     [7:0] sizeBC;                                                         // Size in bytes of beats
logic     [7:0] sizeMask;                                                       // Mask based on size
logic           algnMiss;                                                       // Misaligned to size flag
logic     [2:0] aBeats;                                                         // Number of beats when aligned
logic     [8:0] tBeats;                                                         // Total number of beats (and width adjusted)
logic     [7:0] flitSkip;                                                       // Flits skipped due to mis-aligned address (when beat > flit) 
logic     [7:0] fBCMask;                                                        // Mask based on flit width
logic     [7:0] flitOff;                                                        // Offset within the flit of the first beat in units of beat
logic    [11:0] lenMask;                                                        // Mask based on total length (WRAP only)
logic    [11:0] wrapTo;                                                         // Address we WRAP to
logic    [11:0] wrapFrom;                                                       // Address we WRAP from
logic           wrapAdd;                                                        // Set when WRAP will add a flit
logic     [3:0] flitShift;                                                      // Shift to multiply or divide by "beats per flit"
logic     [5:0] flitsPerBeat;                                                   // Flits in a normal beat
logic     [5:0] flitFirstLoop;                                                  // Flits in first loop
logic     [5:0] flitPerLoop;                                                    // Flits per loop after first loop
logic     [8:0] flitLoops;                                                      // Number of flit loops
logic    [31:0] rregdata;
logic     [1:0] rregmode;
logic     [1:0] rregmode_nxt;
logic     [0:0] rregmode_en;
// ========================================================================//
// Parameter Declarations
// ========================================================================//
// ========================================================================//
// Process parameters and create local derived variables
// ========================================================================//
// ========================================================================//
// Define module I/O
// ========================================================================//
// ============================================
// Clocks and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Forward Channel 0 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_rtr0_nulltgt_f0pipe f0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f0_activity),                                                   // i:1
  .src_req(f0_req),                                                             // i:1
  .src_sop(f0_sop),                                                             // i:1
  .src_eop(f0_eop),                                                             // i:1
  .src_flitdata(f0_flitdata),                                                   // i:36
  .src_ready(f0_ready),                                                         // o:1
  .dst_activity(if0_activity),                                                  // o:1
  .dst_req(if0_req),                                                            // o:1
  .dst_sop(if0_sop),                                                            // o:1
  .dst_eop(if0_eop),                                                            // o:1
  .dst_flitdata(if0_flitdata),                                                  // o:36
  .dst_ready(if0_ready)                                                         // i:1
);
// ============================================
// Forward Channel 1 (LLK manager)
// ============================================
// Forward Channel Pipeline Component
usb4_tc_noc_rtr0_nulltgt_f1pipe f1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(f1_activity),                                                   // i:1
  .src_req(f1_req),                                                             // i:1
  .src_sop(f1_sop),                                                             // i:1
  .src_eop(f1_eop),                                                             // i:1
  .src_flitdata(f1_flitdata),                                                   // i:60
  .src_ready(f1_ready),                                                         // o:1
  .dst_activity(if1_activity),                                                  // o:1
  .dst_req(if1_req),                                                            // o:1
  .dst_sop(if1_sop),                                                            // o:1
  .dst_eop(if1_eop),                                                            // o:1
  .dst_flitdata(if1_flitdata),                                                  // o:60
  .dst_ready(if1_ready)                                                         // i:1
);
// ============================================
// Reverse Channel 0 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_rtr0_nulltgt_r0pipe r0pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir0_activity),                                                  // i:1
  .src_req(ir0_req),                                                            // i:1
  .src_sop(ir0_sop),                                                            // i:1
  .src_eop(ir0_eop),                                                            // i:1
  .src_flitdata(ir0_flitdata),                                                  // i:34
  .src_ready(ir0_ready),                                                        // o:1
  .dst_activity(r0_activity),                                                   // o:1
  .dst_req(r0_req),                                                             // o:1
  .dst_sop(r0_sop),                                                             // o:1
  .dst_eop(r0_eop),                                                             // o:1
  .dst_flitdata(r0_flitdata),                                                   // o:34
  .dst_ready(r0_ready)                                                          // i:1
);
// ============================================
// Reverse Channel 1 (LLK subordinate)
// ============================================
// Reverse Channel Pipeline Component
usb4_tc_noc_rtr0_nulltgt_r1pipe r1pipe (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .src_activity(ir1_activity),                                                  // i:1
  .src_req(ir1_req),                                                            // i:1
  .src_sop(ir1_sop),                                                            // i:1
  .src_eop(ir1_eop),                                                            // i:1
  .src_flitdata(ir1_flitdata),                                                  // i:24
  .src_ready(ir1_ready),                                                        // o:1
  .dst_activity(r1_activity),                                                   // o:1
  .dst_req(r1_req),                                                             // o:1
  .dst_sop(r1_sop),                                                             // o:1
  .dst_eop(r1_eop),                                                             // o:1
  .dst_flitdata(r1_flitdata),                                                   // o:24
  .dst_ready(r1_ready)                                                          // i:1
);
// =======================================================================
// Signal declarations
// =======================================================================
// Write Response Header Fields
// Write Command + Data Sequencer Signals
// Write Command extra packet fields
// Read Data + Status Header fields
// Read Command Sequencer Signals
assign frst_n = rst_n;
// Write Command + Data Sequencer states
parameter S_WCD_HDR = 2'd0;
parameter S_WCD_WD = 2'd1;
parameter S_WCD_WS = 2'd2;
// Read Command + Data + Status Sequencer states
parameter S_RC_HDR = 2'd0;
parameter S_RDS_HDR = 2'd1;
parameter S_RDS_PLD = 2'd2;
// ============================================
// Clock Gating Logic
// ============================================
assign wclkEn = if0_activity || (wcd_state != S_WCD_HDR) || (|wc_cnt);
usb4_tc_noc_rtr0_nulltgt_wcg wcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(wclkEn),                                                               // i:1
  .clkOut(wclk),                                                                // o:1
  .isActive()                                                                   // o:1
);
assign rclkEn = if1_activity || (|rc_cnt) || (|rds_cnt)|| (rds_state != S_RC_HDR);
usb4_tc_noc_rtr0_nulltgt_rcg rcg (
  .clk(clk),                                                                    // i:1
  .rst_n(rst_n),                                                                // i:1
  .enbIn(rclkEn),                                                               // i:1
  .clkOut(rclk),                                                                // o:1
  .isActive()                                                                   // o:1
);
// =======================================================================
// Write Command + Data Path Processing
// =======================================================================
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign wc_bus[35:0] = wc_buf[0];
assign wc_bus[71:36] = ((wcd_state == S_WCD_HDR) && (wc_cnt == 1'd1)) ? if0_flitdata : wc_buf[1];
// ============================================
// Write command flit count
// ============================================
always_ff @(posedge wclk, negedge frst_n)
begin
  if (!frst_n)
    wc_cnt <= #1ps 1'd0;
  else if (wc_cnt_en)
    wc_cnt <= #1ps wc_cnt_nxt;
end

// Flop the ingress port index
always_ff @(posedge wclk, negedge frst_n)
begin
  if (!frst_n)
    wr_portIdx <= #1ps 1'd0;
  else if (wr_portIdx_en)
    wr_portIdx <= #1ps wr_portIdx_nxt;
end

assign r1_dstIdx = wr_portIdx_nxt;
// ============================================
// Write status flit count
// ============================================
always_ff @(posedge wclk, negedge frst_n)
begin
  if (!frst_n)
    ws_cnt <= #1ps 1'd0;
  else if (ws_cnt_en)
    ws_cnt <= #1ps ws_cnt_nxt;
end

always_ff @(posedge wclk, negedge frst_n)
begin
  if (!frst_n)
    wcd_state <= #1ps S_WCD_HDR;
  else if (wcd_state_en)
    wcd_state <= #1ps wcd_state_nxt;
end

always_ff @(posedge wclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      wc_buf[0] <= #1ps {36{1'b0}};
      wc_buf[1] <= #1ps {36{1'b0}};
    end
  else
    begin
      if (wc_buf_en[0])
        wc_buf[0] <= #1ps if0_flitdata;
      if (wc_buf_en[1])
        wc_buf[1] <= #1ps if0_flitdata;
    end
end

assign wc_buf_en = wc_buf_we << wc_cnt;
always_ff @(posedge wclk, negedge frst_n)
begin
  if (!frst_n)
    wregdata <= #1ps {36{1'b0}};
  else if (wregdata_en)
    wregdata <= #1ps wregdata_nxt;
end

always_ff @(posedge wclk, negedge frst_n)
begin
  if (!frst_n)
    wregmode <= #1ps 2'd0;
  else if (wregmode_en)
    wregmode <= #1ps wregmode_nxt;
end

assign writeAddr = wc_bus[54:23];
assign regWAddr = writeAddr[11:2];
assign segIdx = regWAddr[0:0] & 1'd0;
assign flitSeg[0] = if0_flitdata[35:0];
assign regWData = wregdata[31:0];
assign regWEn = wregdata[35:32];
always_comb
begin
  // Defaults
  wcd_state_nxt    = wcd_state;
  wc_cnt_nxt       = wc_cnt;
  ws_cnt_nxt       = ws_cnt;
  if0_ready        = 1'b1;
  ir1_activity     = 1'b0;
  ir1_req          = 1'b0;
  ir1_sop          = 1'b0;
  ir1_eop          = 1'b0;
  wr_portIdx_nxt   = wr_portIdx;
  // Write enables
  wcd_state_en     = 1'b0;
  wc_buf_we        = 1'b0;
  wc_cnt_en        = 1'b0;
  ws_cnt_en        = 1'b0;
  wr_portIdx_en    = 1'b0;
  wregdata_nxt     = wregdata;
  wregdata_en      = 1'b0;
  wregmode_nxt     = wregmode;
  wregmode_en      = 1'b0;
  regWReq          = 1'b0;
  case (wcd_state)
    S_WCD_HDR:
      begin
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if0_req)
          begin
            wc_buf_we     = 1'b1;
            wc_cnt_en     = 1'b1;
            // Check for first flit and record source port
            if( wc_cnt == 1'd0 )
              begin
                wr_portIdx_en  = 1'b1;
                wr_portIdx_nxt = f0_srcIdx;
              end
            // Header transmission is complete
            if (wc_cnt == 1'd1)
              begin
                wcd_state_nxt = S_WCD_WD;
                wcd_state_en  = 1'b1;
                wc_cnt_nxt    = 1'd0;
                wregmode_en   = 1'b1;
                if( writeAddr[32-1:12] == 20'd128 &&  writeAddr[1:0] == 2'd0 && wc_bus[22:20] == 3'd4 && int_awdid == 3'd0 )
                    wregmode_nxt = 2'd1;
                else
                    wregmode_nxt = 2'd0;
              end
            // Continuing header transmission
            else
              wc_cnt_nxt = wc_cnt + 1'd1;
          end
      end
   S_WCD_WD:
      begin
        if (if0_req)
          begin
            if( wregmode == 2'd1 )
              begin
                wregmode_en  = 1'b1;
                wregmode_nxt = 2'd2;
                wregdata_en  = 1'b1;
                wregdata_nxt = flitSeg[segIdx];
              end
            if ( if0_eop)
              begin
                wcd_state_nxt     = S_WCD_WS;
                wcd_state_en      = 1'b1;
                ws_cnt_nxt        = 1'd0;
                ws_cnt_en         = 1'b1;
                ir1_activity      = 1'b1;
              end
          end
      end
    S_WCD_WS:
      begin
        if0_ready    = 1'b0;
        ir1_activity = 1'b1;
        ir1_req      = 1'b1;
        ir1_sop      = (ws_cnt == 1'd0);
        ir1_eop      = (ws_cnt == 1'd0);
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir1_ready)
          begin
            // Header transmission is complete
            if (ws_cnt == 1'd0)
              begin
                ws_cnt_nxt  = 1'd0;
                ws_cnt_en   = 1'b1;
                wcd_state_nxt = S_WCD_HDR;
                wcd_state_en  = 1'b1;
                if( wregmode != 2'd0 )
                  begin
                      regWReq      = 1'b1;
                      wregmode_en  = 1'b1;
                      wregmode_nxt = 2'd0;
                  end
              end
            else
              begin
                ws_cnt_nxt  = ws_cnt + 1'd1;
                ws_cnt_en   = 1'b1;
              end
          end
      end
  endcase
end

// ============================================
// Write Response header field assignments
// ============================================
// Write Command + Data Signal Unpacking
assign int_awqos = wc_bus[3:0];
assign int_awsid = wc_bus[17:15];
assign int_awdid = wc_bus[6:4];
assign int_awid = wc_bus[19:18];
assign int_awbar = 2'd0;
always_comb
begin
  // Set default header to all 0s
  ws_hdr            = {24{1'b0}};
  // Assign over the various fields
  ws_hdr[3:0]  = int_awqos;                                                     // loopback QoS from write command
  ws_hdr[6:4]  = int_awsid;                                                     // loopback SID from write command to DID
  ws_hdr[7]  = 1'b1;                                                            // SoT: not supporting fragmentation yet
  ws_hdr[8]  = 1'b1;                                                            // EoT: not supporting fragmentation yet
  ws_hdr[14:9]  = 6'd3;                                                         // Write response command
  ws_hdr[17:15]  = int_awdid;                                                   // loopback DID from wrtie command to SID
  ws_hdr[23:20] = (wregmode!=2'd0) ? 4'd0 : 4'd3;                               // Success or Address error based on register access mode
  ws_hdr[19:18]   = int_awid;
end

// ============================================
// Generate the flit data for the R1 LLK interface
// ============================================
always_comb
begin
  case(ws_cnt)
    1'd0: ir1_flitdata = ws_hdr[23:0];
    default: ir1_flitdata = {24{1'b0}};
  endcase
end

// =======================================================================
// Read Path Processing
// =======================================================================
// =======================================================================
// Read Command Path Processing
// =======================================================================
// Create incoming wc.bus (may be combinatorial or part flops, part comb)
// This is intended to bypass the buffer for the current packing index
assign rc_bus[59:0] = ((rds_state == S_RC_HDR) && (rc_cnt == 1'd0)) ? if1_flitdata : rc_buf[0];
always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    rc_cnt <= #1ps 1'd0;
  else if (rc_cnt_en)
    rc_cnt <= #1ps rc_cnt_nxt;
end

always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    begin
      rc_buf[0] <= #1ps {60{1'b0}};
    end
  else
    begin
      if (rc_buf_en[0])
        rc_buf[0] <= #1ps if1_flitdata;
    end
end

assign rc_buf_en = rc_buf_we << rc_cnt;
// Flop the ingress port index
always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    rc_portIdx <= #1ps 1'd0;
  else if (rc_portIdx_en)
    rc_portIdx <= #1ps rc_portIdx_nxt;
end

assign r0_dstIdx = rc_portIdx_nxt;
assign int_arIsCMO = 1'b0;
assign int_rplen = (int_arIsCMO) ? 3'd1 : rc_bus[22:20];
assign int_araddr = rc_bus[54:23];
assign int_ardid = rc_bus[6:4];
assign isNarrow = int_arsize < 4'd2;
// ============================================
// Read Data + Status Header field assignments
// ============================================
always_comb
begin
  // Set default header to all 0s
  rds_hdr            = {68{1'b0}};
  // Assign over the various fields
  rds_hdr[3:0]  = rc_bus[3:0];                                                  // loopback QoS from write command
  rds_hdr[6:4]  = rc_bus[17:15];                                                // loopback SID from write command to DID
  rds_hdr[7]  = 1'b1;                                                           // SoT: not supporting fragmentation yet
  rds_hdr[8]  = 1'b1;                                                           // EoT: not supporting fragmentation yet
  rds_hdr[14:9]  = 6'd1;                                                        // Read data / status
  rds_hdr[17:15]  = rc_bus[6:4];                                                // loopback DID from write command to SID
  rds_hdr[19:18]   = rc_bus[19:18];                                             // loopback transaction id
  rds_hdr[22:20] = int_rplen;
  rds_hdr[30:23]  = (int_arburst==2'd2) ?  8'(int_araddr>>int_arsize[2:0]) : int_araddr[7:0];
  rds_hdr[33:31]  = int_arsize[2:0];
  rds_hdr[35:34] = int_arburst;
end

// ============================================
// Read Command + Data + Status flit sequencer
// ============================================
always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    rds_cnt <= #1ps 1'd0;
  else if (rds_cnt_en)
    rds_cnt <= #1ps rds_cnt_nxt;
end

always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    rds_state <= #1ps S_RC_HDR;
  else if (rds_state_en)
    rds_state <= #1ps rds_state_nxt;
end

always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    oLoop <= #1ps 9'd0;
  else if (oLoop_en)
    oLoop <= #1ps oLoop_nxt;
end

always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    iLoop <= #1ps 6'd0;
  else if (iLoop_en)
    iLoop <= #1ps iLoop_nxt;
end

assign int_arsize = 4'(rc_bus[57:55]);
assign int_arburst = rc_bus[59:58];
assign tmp_arsize = ({{9{1'b0}},int_rplen} == 12'd1) ? 4'd0 : int_arsize;
assign sizeBC = 8'd1<<tmp_arsize;                                               // Size in bytes of beats
assign sizeMask = sizeBC - 8'd1;                                                // Mask based on size
assign algnMiss = ({{5{1'b0}},int_rplen} & sizeMask) != 8'd0;                   // Misaligned to size flag
assign aBeats = int_rplen>>tmp_arsize;                                          // Number of beats when aligned
assign tBeats = {{6{1'b0}},aBeats} + {{8{1'b0}},algnMiss};                      // Total number of beats (and width adjusted)
assign flitSkip = (int_araddr[7:0] & sizeMask) >> 4'd2;                         // Flits skipped due to mis-aligned address (when beat > flit) 
assign fBCMask = 8'd3;                                                          // Mask based on flit width
assign flitOff = (int_araddr[7:0] & fBCMask) >> tmp_arsize;                     // Offset within the flit of the first beat in units of beat
assign lenMask = ({{9{1'b0}},int_rplen} - 12'd1);                               // Mask based on total length (WRAP only)
assign wrapTo = (int_araddr[11:0] & ~lenMask);                                  // Address we WRAP to
assign wrapFrom = wrapTo + {{9{1'b0}},int_rplen};                               // Address we WRAP from
assign wrapAdd = (wrapTo!=int_araddr[11:0]) && ((wrapFrom[7:0]&fBCMask) != 8'd0);// Set when WRAP will add a flit
assign flitsPerBeat = 6'b1 << flitShift;                                        // Flits in a normal beat
always_comb
begin
  if( tmp_arsize >= 4'd2 )
    begin
      // Since size can be more than 1 flit, the offset within the flit can affect the flit count
      flitShift    = tmp_arsize - 4'd2;
      flitLoops    = tBeats;
      if( int_arburst == 2'd0 )                                                 // FIXED
        begin
          flitFirstLoop = flitsPerBeat - flitSkip[5:0];
          flitPerLoop   = flitsPerBeat - flitSkip[5:0];
        end
      else if( int_arburst == 2'd2 )                                            // WRAP
        begin
          flitFirstLoop = flitsPerBeat;
          flitPerLoop   = flitsPerBeat;
        end
      else
        begin
          flitFirstLoop = flitsPerBeat - flitSkip[5:0];
          flitPerLoop   = flitsPerBeat;
        end
    end
  else
    begin
      // Since size is less than 1 flit, the size offset alone determines the flit count
      flitShift     = 4'd2 - tmp_arsize;
      flitPerLoop   = 6'd1;
      flitFirstLoop = 6'd1;
      if( isNarrow || int_arburst == 2'd0 )                                     // Narrow Read or FIXED
          flitLoops = tBeats;
      else if( int_arburst == 2'd2 )                                            // WRAP
        begin
          flitLoops = 9'(({{5{1'b0}},tBeats} + {{6{1'b0}},flitOff} + (14'd1<<flitShift) - 14'd1) >> flitShift) + {{8{1'b0}},wrapAdd};
        end
      else
        begin
          flitLoops = 9'(({{5{1'b0}},tBeats} + {{6{1'b0}},flitOff} + (14'd1<<flitShift) - 14'd1) >> flitShift);
        end
    end
end

always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    rregdata <= #1ps 32'd0;
  else if (regRReq)
    rregdata <= #1ps regRData;
end

always_ff @(posedge rclk, negedge frst_n)
begin
  if (!frst_n)
    rregmode <= #1ps 2'd0;
  else if (rregmode_en)
    rregmode <= #1ps rregmode_nxt;
end

assign regRAddr = int_araddr[11:2];
always_comb
begin
  // Defaults
  rds_state_nxt = rds_state;
  rds_cnt_nxt   = rds_cnt;
  rc_cnt_nxt    = rc_cnt;
  ir0_activity  = 1'b0;
  ir0_req       = 1'b0;
  ir0_sop       = 1'b0;
  ir0_eop       = 1'b0;
  ir0_flitdata  = {34{1'b0}};
  rc_portIdx_nxt = rc_portIdx;
  // Write enables
  rds_state_en  = 1'b0;
  rds_cnt_en    = 1'b0;
  rc_cnt_en     = 1'b0;
  rc_buf_we     = 1'b0;
  rc_portIdx_en = 1'b0;
  iLoop_nxt     = iLoop;
  iLoop_en      = 1'b0;
  oLoop_nxt     = oLoop;
  oLoop_en      = 1'b0;
  if1_ready     = 1'b0;
  rregmode_nxt     = rregmode;
  rregmode_en      = 1'b0;
  regRReq          = 1'b0;
  case (rds_state)
    S_RC_HDR:
      begin
        if1_ready = 1'b1;
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (if1_req)
          begin
            rc_buf_we     = 1'b1;
            rc_cnt_en     = 1'b1;
            // Check for first flit and record source port
            if( rc_cnt == 1'd0 )
              begin
                rc_portIdx_en  = 1'b1;
                rc_portIdx_nxt = f1_srcIdx;
              end
            // Header reception is complete
            if (rc_cnt == 1'd0)
              begin
                rds_state_nxt = S_RDS_HDR;
                rds_state_en  = 1'b1;
                rc_cnt_nxt    = 1'd0;
                ir0_activity  = 1'b1;
                rregmode_en   = 1'b1;
                if( int_araddr[32-1:12] == 20'd128 && int_araddr[1:0] == 2'd0 && int_rplen == 3'd4 && int_ardid == 3'd0 )
                  begin
                    regRReq      = 1'b1;
                    rregmode_nxt = 2'd1;
                  end
                else
                    rregmode_nxt = 2'd0;
              end
            // Continuing header reception
            else
              rc_cnt_nxt = rc_cnt + 1'd1;
          end
      end
    S_RDS_HDR:
      begin
        ir0_activity  = 1'b1;
        ir0_req   = 1'b1;
        ir0_sop   = (rds_cnt == 1'd0);
        case(rds_cnt)
          1'd0: ir0_flitdata = rds_hdr[33:0];
          1'd1: ir0_flitdata = rds_hdr[67:34];
          default: ir0_flitdata = {34{1'b0}};
        endcase
        // Update the header fragment count and generate the ready back to the ingress pipe stage
        if (ir0_ready)
          begin
            // Header transmission is complete
            if (rds_cnt == 1'd1)
              begin
                rds_cnt_nxt      = 1'd0;
                rds_cnt_en       = 1'b1;
                rds_state_nxt    = S_RDS_PLD;
                rds_state_en     = 1'b1;
                oLoop_en         = 1'b1;
                oLoop_nxt        = flitLoops;
                iLoop_en         = 1'b1;
                iLoop_nxt        = flitFirstLoop;
              end
            // Continuing header transmission
            else
              begin
                rds_cnt_nxt = rds_cnt + 1'd1;
                rds_cnt_en  = 1'b1;
              end
          end
      end
   S_RDS_PLD:
      begin
        ir0_activity  = 1'b1;
        ir0_req       = 1'b1;
        ir0_eop       = oLoop==9'd1 && iLoop==6'd1;
        if( rregmode == 2'd1 )
            ir0_flitdata = {1{ 2'b0, rregdata[31:0] }};
        else
          begin
            ir0_flitdata  = {1{2'b11,32'd0}};
          end
        if (ir0_ready)
          begin
          if( rregmode == 2'd1 )
            begin
              rregmode_en  = 1'b1;
              rregmode_nxt = 2'd2;
            end
          if( rregmode == 2'd2 )
            begin
              rregmode_en  = 1'b1;
              rregmode_nxt = 2'd3;
            end
            if (ir0_eop)
              begin
                rds_state_nxt = S_RC_HDR;
                rds_state_en  = 1'b1;
              end
            else
              begin
                iLoop_en = 1'b1;
                if( iLoop==6'd1 )
                  begin
                    iLoop_nxt = flitPerLoop;
                    oLoop_en  = 1'b1;
                    oLoop_nxt = oLoop - 9'd1;
                  end
                else
                  iLoop_nxt = iLoop - 6'd1;
              end
          end
      end
  endcase
end

endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_f0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [35:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [35:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_nulltgt_f0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:36
  .dst_flitdata(dst_flitdata)                                                   // o:36
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_f0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [35:0] src_flitdata,
  output logic    [35:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_f1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [59:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [59:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_nulltgt_f1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:60
  .dst_flitdata(dst_flitdata)                                                   // o:60
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_f1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [59:0] src_flitdata,
  output logic    [59:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_r0pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [33:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [33:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_nulltgt_r0pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:34
  .dst_flitdata(dst_flitdata)                                                   // o:34
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_r0pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [33:0] src_flitdata,
  output logic    [33:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_r1pipe (
  input  wire            clk,
  input  wire            rst_n,
  // src
  input  wire            src_activity,                                          // Upcoming activity indicator
  input  wire            src_req,                                               // Flit transfer request
  input  wire            src_sop,                                               // Start of packet indicator
  input  wire            src_eop,                                               // End of packet indicator
  input  wire     [23:0] src_flitdata,                                          // Flit data
  output logic           src_ready,                                             // Flit transfer ready
  // dst
  output logic           dst_activity,                                          // Upcoming activity indicator
  output logic           dst_req,                                               // Flit transfer request
  output logic           dst_sop,                                               // Start of packet indicator
  output logic           dst_eop,                                               // End of packet indicator
  output logic    [23:0] dst_flitdata,                                          // Flit data
  input  wire            dst_ready                                              // Flit transfer ready
);

logic           frst_n;
// ============================================
// Clock and reset
// ============================================
// ============================================
// Test Mode + Clock Gating Override
// ============================================
// ============================================
// Source Port (LLK subordinate)
// ============================================
// ============================================
// Destination Port (LLK manager)
// ============================================
// ============================================
// Half reset synchronizer
// ============================================
assign frst_n = rst_n;
// ===========================================
// Channel FIFO
// ===========================================
usb4_tc_noc_rtr0_nulltgt_r1pipe_cfifo cfifo (
  .clk(clk),                                                                    // i:1
  .rst_n(frst_n),                                                               // i:1
  .wreq(src_req),                                                               // i:1
  .wact(src_activity),                                                          // i:1
  .ract(dst_activity),                                                          // o:1
  .wrdy(src_ready),                                                             // o:1
  .rreq(dst_ready),                                                             // i:1
  .rrdy(dst_req),                                                               // o:1
  .src_sop(src_sop),                                                            // i:1
  .dst_sop(dst_sop),                                                            // o:1
  .src_eop(src_eop),                                                            // i:1
  .dst_eop(dst_eop),                                                            // o:1
  .src_flitdata(src_flitdata),                                                  // i:24
  .dst_flitdata(dst_flitdata)                                                   // o:24
);
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_r1pipe_cfifo (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            wreq,
  input  wire            wact,
  output logic           ract,
  output logic           wrdy,
  input  wire            rreq,
  output logic           rrdy,
  input  wire            src_sop,
  output logic           dst_sop,
  input  wire            src_eop,
  output logic           dst_eop,
  input  wire     [23:0] src_flitdata,
  output logic    [23:0] dst_flitdata
);

logic     [0:0] crun;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    crun <= #1ps 1'd0;
  else
    crun <= #1ps ract;
end

assign wrdy = rreq && crun;
assign rrdy = wreq && crun;
assign ract = wreq || wact;
assign dst_sop = src_sop;
assign dst_eop = src_eop;
assign dst_flitdata = src_flitdata;
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_wcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

// Copyright (c) 2013-2025 by Cadence Design Systems Inc.  ALL RIGHTS RESERVED.
// These coded instructions, statements, and computer programs are the copyrighted
// works and confidential proprietary information of Cadence Design Systems Inc.
// They may not be modified, copied, reproduced, distributed, or disclosed to
// third parties in any manner, medium, or form, in whole or in part, without the
// prior written consent of Cadence Design Systems Inc.

module usb4_tc_noc_rtr0_nulltgt_rcg (
  input  wire            clk,
  input  wire            rst_n,
  input  wire            enbIn,                                                 // Enable input signal
  output wire            clkOut,                                                // Output clock
  output wire            isActive                                               // Output activity signal
);

logic     [0:0] holdEnable;
always_ff @(posedge clk, negedge rst_n)
begin
  if (!rst_n)
    holdEnable <= #1ps 1'b1;
  else
    holdEnable <= #1ps enbIn;
end

assign isActive = holdEnable;
usb4_tc_noc_xtgated_clock midlevel_cg (
  .xtout(clkOut),                                                               // (external)
  .xten(isActive),                                                              // (external)
  .xtclk(clk)                                                                   // (external)
);
// Make sure our standard primitives are copied over
endmodule

