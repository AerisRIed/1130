`include "cdn_u4_usb4_test_base.sv"

`ifdef DENALI_USB4_VIP
`include "cdn_u4_usb4_vip_test_base.sv"
`endif
