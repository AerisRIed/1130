`include"cdn_u4_dp_base_sequence.sv"
`include"cdn_u4_dp_virtual_sequence.sv"
`include"cdn_u4_dp_start_up_sequence.sv"

