`include"usb4_base_sequence.sv"
//`include"usb4_cl1_entry_device_request_sequence.sv"
//`include"usb4_cl1_entry_host_request_sequence.sv"
//`include"usb4_cl1_exit_host_request_sequence.sv"
