`include "passive_master_usb4_tc_noc_cmn_cdb_config.sv"
`include "active_slave_usb4_tc_noc_cmn_cdb_config.sv"
`include "passive_master_usb4_tc_noc_tc_reg_config.sv"
`include "active_slave_usb4_tc_noc_tc_reg_config.sv"
`include "passive_master_usb4_tc_noc_usb_sub_sys_config.sv"
`include "active_slave_usb4_tc_noc_usb_sub_sys_config.sv"
`include "passive_master_usb4_tc_noc_pam3_sub_sys_config.sv"
`include "active_slave_usb4_tc_noc_pam3_sub_sys_config.sv"
`include "passive_master_usb4_tc_noc_apb_tgt_config.sv"
`include "active_slave_usb4_tc_noc_apb_tgt_config.sv"
`include "passive_master_usb4_tc_noc_xcvr_ln_0_config.sv"
`include "active_slave_usb4_tc_noc_xcvr_ln_0_config.sv"
`include "passive_slave_usb4_tc_noc_apb_mstr_config.sv"
`include "active_master_usb4_tc_noc_apb_mstr_config.sv"
`include "passive_slave_usb4_tc_noc_cdb_config.sv"
`include "active_master_usb4_tc_noc_cdb_config.sv"
