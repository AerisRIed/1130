`include "cdn_usb_phy_reg_seq.sv"
