//package cdn_phy_params;

parameter DATA_WIDTH = 32; //TBD

parameter POWER_IDLE = 6'b00_0000;
parameter POWER_A0   = 6'b00_0001;
parameter POWER_A1   = 6'b00_0010;
parameter POWER_A2   = 6'b00_0100;
parameter POWER_A3   = 6'b00_1000;
parameter POWER_A4   = 6'b01_0000;
parameter POWER_A5   = 6'b10_0000;

//endpackage

//import cdn_phy_params::*;
