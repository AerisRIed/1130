`define PAIR_OFFSET		12'h200

`define PHY_RX_MRGN_CTRL_0	12'h000 + `PAIR_OFFSET
`define PHY_RX_MRGN_CTRL_1	12'h001 + `PAIR_OFFSET
`define PHY_EL_BUF_CTRL		12'h002 + `PAIR_OFFSET
`define PHY_RX_CTRL_0		12'h003 + `PAIR_OFFSET
`define PHY_RX_CTRL_1		12'h004 + `PAIR_OFFSET
`define PHY_RX_CTRL_2		12'h005 + `PAIR_OFFSET
`define PHY_RX_CTRL_3		12'h006 + `PAIR_OFFSET
`define PHY_EL_BUF_LOC_UP_FRQ	12'h007 + `PAIR_OFFSET
`define PHY_RX_CTRL_4		12'h008 + `PAIR_OFFSET
`define PHY_RX_CTRL_5		12'h009 + `PAIR_OFFSET

`define PHY_TX_CTRL_0		12'h400 + `PAIR_OFFSET
`define PHY_TX_CTRL_1		12'h401 + `PAIR_OFFSET
`define PHY_TX_CTRL_2		12'h402 + `PAIR_OFFSET
`define PHY_TX_CTRL_3		12'h403 + `PAIR_OFFSET
`define PHY_TX_CTRL_4		12'h404 + `PAIR_OFFSET
`define PHY_TX_CTRL_5		12'h405 + `PAIR_OFFSET
`define PHY_TX_CTRL_6		12'h406 + `PAIR_OFFSET
`define PHY_TX_CTRL_7		12'h407 + `PAIR_OFFSET
`define PHY_TX_CTRL_8		12'h408 + `PAIR_OFFSET
`define PHY_TX_CTRL_9		12'h409 + `PAIR_OFFSET

`define PHY_CMN_CTRL_0       	12'h800 + `PAIR_OFFSET
`define PHY_NEL_CTRL_0       	12'h801 + `PAIR_OFFSET
