`include "cdn_usb_phy_reg_try_test.sv"
`include "cdn_usb_phy_illegal_address_reg_test.sv"
