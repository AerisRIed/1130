`ifndef VALUE_DEFINES__SVH
`define VALUE_DEFINES__SVH
//NOTE:just a demo from torrent
    // `define PHY_PIPE_CMN_CTRL            16'hC000
    // `define PHY_PIPE_COM_LOCK_CFG1       16'hC002
    // `define PHY_PIPE_COM_LOCK_CFG2       16'hC003
    // `define PHY_PIPE_SYNC_LOCK_CFG       16'hC004
    // `define PHY_PIPE_RCV_DET_INH         16'hC006
    // `define PHY_PIPE_RX_ELEC_IDLE_DLY    16'hC007
    // `define PHY_ISO_CMN_CTRL1            16'hC008
    // `define PHY_ISO_CMN_CTRL2            16'hC009
    // `define PHY_ISO_CMN_CTRL3            16'hC00A
    // `define PHY_STATE_CHG_TIMEOUT        16'hC00C
    // `define DTB_DATA_LOW                 16'hC00D
    // `define DTB_DATA_HIGH                16'hC00E
    // `define PHY_AUTO_CFG_SPDUP           16'hC00F
    // `define PHY_PMA_LANE_MAP             16'hC010
    // `define PHY_LANE_OFF_CTL             16'hC011
    // `define PHY_USB_INTERRUPT_STS        16'hC014
    // `define PHY_DP_INTERRUPT_STS         16'hC015
    // `define PHY_PIPE_USB3_GEN2_PRE_CFG0  16'hC018
    // `define PHY_PIPE_USB3_GEN2_PRE_CFG1  16'hC019
    // `define PHY_PIPE_USB3_GEN2_POST_CFG0 16'hC01A
    // `define PHY_PIPE_USB3_GEN2_POST_CFG1 16'hC01B

    // `define PHY_USB3_ISO_TX_CTRL         16'hD000
    // `define PHY_USB3_ISO_TX_FSLF         16'hD005
    // `define PHY_USB3_ISO_TX_DATA_LO      16'hD006
    // `define PHY_USB3_ISO_TX_DATA_HI      16'hD007
    // `define PHY_USB3_ISO_RX_CTRL         16'hD008
    // `define PHY_USB3_USB_BER_CNT         16'hD00C
    // `define PHY_USB3_ISO_RX_DATA_LO      16'hD00E
    // `define PHY_USB3_ISO_RX_DATA_HI      16'hD00F
    // `define PHY_DP_ISO_TC_CTRL1          16'hD010
    // `define PHY_DP_ISO_TC_CTRL2          16'hD011

    // `define PHY_PMA_CMN_CTRL1            16'hE000
    // `define PHY_PMA_CMN_CTRL2            16'hE001
    // `define PHY_PMA_SSM_STATE            16'hE002
    // `define PHY_PMA_PLL_CTRL             16'hE003
    // `define PHY_PMA_ISO_CMN_CTRL         16'hE004
    // `define PHY_PMA_ISO_PLL_CTRL0        16'hE005
    // `define PHY_PMA_ISO_PLL_CTRL1        16'hE006
    // `define PHY_PMA_PLL0_SM_STATE        16'hE00B
    // `define PHY_PMA_PLL1_SM_STATE        16'hE00C
    // `define PHY_PMA_ISOLATION_CTRL       16'hE00F

    // `define PHY_PMA_XCVR_CTRL            16'hF000
    // `define PHY_PMA_XCVR_LPBK            16'hF001
    // `define PHY_PMA_PI_POS               16'hF002
    // `define PHY_PMA_ISO_XCVR_CTRL        16'hF003
    // `define PHY_PMA_ISO_TX_LPC_LO        16'hF004
    // `define PHY_PMA_ISO_TX_LPC_HI        16'hF005
    // `define PHY_PMA_ISO_TX_DMPH_LO       16'hF006
    // `define PHY_PMA_ISO_TX_DMPH_HI       16'hF007
    // `define PHY_PMA_ISO_TX_FSLF          16'hF008
    // `define PHY_PMA_ISO_TX_MGN           16'hF009
    // `define PHY_PMA_ISO_LINK_MODE        16'hF00A
    // `define PHY_PMA_ISO_PWRST_CTRL       16'hF00B
    // `define PHY_PMA_ISO_RX_EQ_CTRL       16'hF00D
    // `define PHY_PMA_ISO_RX_DATA_LO       16'hF00E
    // `define PHY_PMA_ISO_RX_DATA_HI       16'hF00F
    // `define PHY_PMA_PSM_STATE_LO         16'hF010
    // `define PHY_PMA_PSM_STATE_HI         16'hF011

    `define TGT_APB_ADDR_WIDTH              32
    `define TGT_APB_DATA_WIDTH              32
`endif