`include"cdn_u4_pcie_test_base.sv"

