/* ------------------------------------------------------------------------------
--
-- CADENCE Copyright (c) 2025
-- Cadence Design Systems, Inc.
-- All rights reserved.
--
-- 
-- This work may not be copied, modified, re-published, uploaded, executed, or
-- distributed in any way, in any medium, whether in whole or in part, without
-- prior written permission from Cadence Design Systems, Inc.
--------------------------------------------------------------------------------- */


class dut_usb4_tc_noc_env_vip_container extends uvm_env;

   // pointer to the env configuration
   dut_usb4_tc_noc_env_cfg env_cfg;

   // reference to the routing model
   cdn_stg_routing_model routing_model;

   // configure this string from above to set the path to the module where the VIP
   // wrapper modules are instantiated
   string vip_wrapper_modules_path;

   cdn_stg_apb_basic_env_port cmn_cdb;
   cdn_stg_apb_basic_env_port tc_reg;
   cdn_stg_apb_basic_env_port usb_sub_sys;
   cdn_stg_apb_basic_env_port pam3_sub_sys;
   cdn_stg_apb_basic_env_port apb_tgt;
   cdn_stg_apb_basic_env_port xcvr_ln_0;


   cdn_stg_apb_basic_env_port apb_mstr;
   cdn_stg_apb_basic_env_port cdb;


   `uvm_component_utils_begin(dut_usb4_tc_noc_env_vip_container)
	`uvm_field_string(vip_wrapper_modules_path, UVM_ALL_ON)
   `uvm_component_utils_end


   function new(string name="dut_usb4_tc_noc_env_vip_container", uvm_component parent=null);
	super.new(name,parent);
   endfunction

   extern virtual function void apb_build_code();
   extern virtual function void apb_config_code();

   /*
    *
    * VIP agent instances
    *
    */

   /*
    *
    * build_phase
    *
    */
   virtual function void build_phase(uvm_phase phase);
	super.build_phase(phase);

	// code generated by the VIP bundles to build the VIP agents
        apb_build_code();
   endfunction


   /*
    *
    * connect_phase
    *
    */
   virtual function void connect_phase(uvm_phase phase);
      	super.connect_phase(phase);

   endfunction


   /*
    *
    * end_of_elaboration_phase
    *
    */
   virtual function void end_of_elaboration_phase(uvm_phase phase);
	super.end_of_elaboration_phase(phase);

	// code generated by the VIP bundles to...
	// configure non-SOMA based features
        apb_config_code();

   endfunction


   /*
    *
    * start_of_simulation_phase
    *
    */
   virtual function void start_of_simulation_phase(uvm_phase phase);
	super.start_of_simulation_phase(phase);

	// configure the memory maps of each VIP agent
	routing_model.configure_all_vip_agents_memory_maps();
   endfunction

endclass

