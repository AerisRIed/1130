extern task write_dp_1p62_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_1p62_none_int_100p0_pll0_None_ssc_pll1_Enable_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_10_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_13p5_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_20_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_2p7_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_5p4_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_8p1_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_2p7_none_int_100p0_pll0_None_ssc_pll1_Enable_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_10_none_int_100p0_pll0_None_ssc_pll1_Enable_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_13p5_none_int_100p0_pll0_None_ssc_pll1_Enable_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_20_none_int_100p0_pll0_None_ssc_pll1_Enable_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_5p4_none_int_100p0_pll0_None_ssc_pll1_Enable_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_dp_8p1_none_int_100p0_pll0_None_ssc_pll1_Enable_ssc_pg_reg(int dp_lane_num, int de_emphasis, int swing, bit flip_flag);
extern task write_usb_tcam_gen1_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen2_none_int_24p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen2_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen1_none_int_100p0_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen1_none_int_19p2_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen1_none_int_19p2_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen1_none_int_24p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen1_none_int_24p0_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen2_none_int_100p0_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen2_none_int_19p2_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen2_none_int_19p2_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb_tcam_gen2_none_int_24p0_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb4_tcam_none_int_100p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb4_tcam_none_int_100p0_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb4_tcam_none_int_19p2_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb4_tcam_none_int_19p2_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb4_tcam_none_int_24p0_pll0_None_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
extern task write_usb4_tcam_none_int_24p0_pll0_Enable_ssc_pll1_None_ssc_pg_reg(int lane_num, string IO_USB_TCAM, bit flip_flag);
