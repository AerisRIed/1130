`include"cdn_u4_usb32_base_sequence.sv"
`include"cdn_u4_usb32_lowpower_base_sequence.sv"
//`include"u32_u1_entry_exit_sequence.sv"
//`include"u32_u2_entry_exit_sequence.sv"
//`include"u32_u3_entry_exit_sequence.sv"

