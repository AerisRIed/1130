// Memory Define Include File
//
// Each of the lines below represents a memory module. When defined, the memory is implemented
// by an external macro. When commented out, the memory is implemented using internal flops.

// `define USB4_TC_NOC_TPRAM_8_35_AWN_RAWS 1
// `define USB4_TC_NOC_TPRAM_8_25_AWN_RAWS 1
// `define USB4_TC_NOC_TPRAM_8_37_AWN_RAWS 1
// `define USB4_TC_NOC_TPRAM_8_61_AWN_RAWS 1
