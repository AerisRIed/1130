  int reg_access_mbx_value;
  bit pending_update = 0;
  bit di_control_write;
  bit try_read_in_progress;
  bit concurrent_reg = 0;
