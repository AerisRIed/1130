`include"usb32_base_sequence.sv"
`include"usb32_u1_entry_device_request_sequence.sv"
`include"usb32_u1_entry_host_request_sequence.sv"
`include"usb32_u1_exit_host_request_sequence.sv"
