/*
 * This empty include file is generated and `included in the compile flow.
 * This allows you to create your own file (of the same name) in your own
 * directory and `include your dut_usb4_tc_noc_tb_test_pkg extensions.
 *
 * Your own files can be included in the compile flow by:
 * 1. create <my extensions dir>/test_pkg/dut_usb4_tc_noc_tb_test_pkg_usr.sv
 *    > `include your own test package extensions files
 * 2. include <my extensions dir>/tb_pkg in the compile flow
 *    > stg -sim ... -irunopts "-incdir <my extensions dir>/test_pkg" ...
 *    or 
 *    > irun ... -incdir <my extensions dir>/test_pkg ...
 *
 */
