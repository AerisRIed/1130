`include"cdn_u4_dp_test_base.sv"


