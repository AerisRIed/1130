`include "cdn_phy_bring_up_seq.sv"