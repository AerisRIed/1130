//-----------------------------------------------------------------------------
//    This confidential and proprietary HDL soft description of a Hardware
//    component may be used only as authorized by a licensing agreement from
//    Cadence. In the event of publication,the following notice 
//    is applicable:
//
//                       (C) COPYRIGHT 2016 Cadence
//                         ALL RIGHTS RESERVED
//
//     The entire notice above must be reproduced on all authorized
//     copies of this code.
//-----------------------------------------------------------------------------
//-----------------------------------------------------------------------------
//
// Filename        : timberwolf_testchip.sv
// Author          : Zhenwei Liu
// Abstract        : This is Testchip module for the Timberwolf 4nm project. It 
//                   contains the following components:
//                        - Testchip pads (TSMC IO, DDR IO, DDR IO Calibration)
//                        - Timberwolf USB Type-C PHY IP (2-lane)
//                        - PAM3 PMA IP (1-lane)
//                        - JTAG TAP controller
//                        - NoC
//                        - Testchip registers
// 
//-----------------------------------------------------------------------------


module timberwolf_testchip (
//--------------------------------------------------
// Supply/Ground Pads
//--------------------------------------------------
`ifdef CDNS_PHY_PWR_AWARE // @RELEASE@
// *******************************
// PHY Power pins
// *******************************
input                           agnd,
input                           avdd_clk,
input                           avdd_h,
input                           avdd,
input                           avdd_tx0,
input                           avdd_tx1,
input                           avdd_tx2,
input                           avdd_tx3,
input                           avdd_rx,
input                           cmn_aonvdd,
input                           vdd,
`endif // @RELEASE@
// *******************************
// PAM3 Power pins
// *******************************
`ifdef CDNS_PMA_PWR_AWARE // @RELEASE@

`endif // @RELEASE@
// *******************************
// Testchip Power pins
// *******************************
`ifdef CDNS_TC_PWR_AWARE // @RELEASE@
input                           gnd,
input                           vdd,
input                           vddio,
input                           vddq,
`endif // @RELEASE@
//--------------------------------------------------
// System Clocks
//--------------------------------------------------
input                           cmn_refclk0_p_phy,
input                           cmn_refclk0_m_phy,
inout                           cmn_refclk1_p_phy,
inout                           cmn_refclk1_m_phy,
input                           cmn_refclk0_p_pam3,
input                           cmn_refclk0_m_pam3,
inout                           cmn_refclk1_p_pam3,
inout                           cmn_refclk1_m_pam3,
input                           cmn_refclk0_int,
input                           cmn_refclk1_int,

//--------------------------------------------------
// NoC Interface
//--------------------------------------------------
input                           noc_clk,
input                           noc_reset_n,

//--------------------------------------------------
// uC clock
//--------------------------------------------------
input                           uc_clk,

//--------------------------------------------------
// TC reset
//--------------------------------------------------
input                           tc_reset_n,

//--------------------------------------------------
// PMA External Interface
// MP PHY Interface
//--------------------------------------------------
//USB Type-C PHY
inout                           xcvr_p_ln_0_phy,
inout                           xcvr_m_ln_0_phy,
inout                           xcvr_p_ln_1_phy,
inout                           xcvr_m_ln_1_phy,
inout                           xcvr_p_ln_2_phy,
inout                           xcvr_m_ln_2_phy,
inout                           xcvr_p_ln_3_phy,
inout                           xcvr_m_ln_3_phy,

input                           cmn_rext_phy,

inout                           atb_0_phy,
inout                           atb_1_phy,
//PAM3 PMA
inout                           xcvr_p_ln_0_pam3,
inout                           xcvr_m_ln_0_pam3,

input                           cmn_rext_pam3,

inout                           atb_0_pam3,
inout                           atb_1_pam3,

output                          test_clk,
input                           iddq_en,

input                           ddr_rext,
//--------------------------------------------------
// TAP Interface
//--------------------------------------------------
input  [1:0]                    sel_tap,
input                           tap_tck,
input                           tap_tms,
input                           tap_trst_n,
input                           tap_tdi,
output                          tap_tdo,

//--------------------------------------------------
// uC debugger TAP Interface
//--------------------------------------------------
input                           uc_tap_tck,
input                           uc_tap_tms,
input                           uc_tap_trst_n,
input                           uc_tap_tdi,
output                          uc_tap_tdo,

//--------------------------------------------------
// AUX/Sideband Interface
//--------------------------------------------------


//--------------------------------------------------
// PCS PIPE external Interface
//--------------------------------------------------
// *******************************
// Common pins
// *******************************
output                          pipe_clk_max,
input                           pipe_reset_n,
input                           pipe_rate,
input                           pipe_clk_max_req,
output                          pipe_clk_max_ack,
input    [2-1:0]                pipe_powerdown,
input                           pipe_pll0_en,
output                          pipe_pll0_ok,
output                          pma_cmn_ready,
output                          phy_interrupt,
input                           typec_conn_dir,
// *******************************
// Lane0 RX pins
// *******************************                        
output                          pipe_l00_rx_clk,
output                          pipe_l00_phy_status,
inout    [32-1:0]               pipe_l00_rx_data,
output   [8-1:0]                pipe_l00_p2m_messagebus,
output                          pipe_l00_rx_start_block,
inout                           pipe_l00_rx_data_valid,
output                          pipe_l00_rx_valid,
output   [3-1:0]                pipe_l00_rx_standby_status,
output                          pipe_l00_rx_elec_idle,
input                           pipe_l00_rx_standby,
input                           pipe_l00_rx_termination,
input                           pipe_l00_rx_eq_training,
// *******************************
// Lane0 TX pins
// *******************************              
input                           pipe_l00_clk,
input    [32-1:0]               pipe_l00_tx_data,
input    [8-1:0]                pipe_l00_m2p_messagebus,
input                           pipe_l00_tx_start_block,
input                           pipe_l00_tx_data_valid,
input                           pipe_l00_tx_det_rx_lpbk,
input                           pipe_l00_tx_elec_idle,
input    [3-1:0]                pipe_l00_powerdown,
input    [2-1:0]                pipe_l00_rate,
// *******************************
// Lane1 RX pins
// *******************************              
output                          pipe_l01_rx_clk,
output                          pipe_l01_phy_status,
inout    [32-1:0]               pipe_l01_rx_data,
output   [8-1:0]                pipe_l01_p2m_messagebus,
output                          pipe_l01_rx_start_block,
inout                           pipe_l01_rx_data_valid,
output                          pipe_l01_rx_valid,
output   [3-1:0]                pipe_l01_rx_standby_status,
output                          pipe_l01_rx_elec_idle,
input                           pipe_l01_rx_standby,
input                           pipe_l01_rx_termination,
input                           pipe_l01_rx_eq_training,
// *******************************
// Lane1 TX pins
// *******************************             
input                           pipe_l01_clk,
input    [32-1:0]               pipe_l01_tx_data,
input    [8-1:0]                pipe_l01_m2p_messagebus,
input                           pipe_l01_tx_start_block,
input                           pipe_l01_tx_data_valid,
input                           pipe_l01_tx_det_rx_lpbk,
input                           pipe_l01_tx_elec_idle,
input    [3-1:0]                pipe_l01_powerdown,
input    [2-1:0]                pipe_l01_rate    
);
 
/****************************************************************************\
|*                                                                          *|
|*      Internal wire/reg Definition                                        *|
|*                                                                          *|
\****************************************************************************/
//--------------------------------------------------
// System Clocks
//--------------------------------------------------
wire                            pad_cmn_refclk0_int;
wire                            pad_cmn_refclk1_int;

//--------------------------------------------------
// NoC Interface
//--------------------------------------------------
wire                            pad_noc_clk;
wire                            pad_noc_reset_n;

//--------------------------------------------------
// uC clock
//--------------------------------------------------
wire                            pad_uc_clk;

//--------------------------------------------------
// TC reset
//--------------------------------------------------
wire                            pad_tc_reset_n;

//--------------------------------------------------
// PMA External Interface
// MP PHY Interface
//--------------------------------------------------
wire                            pad_test_clk;
wire                            pad_iddq_en;

//--------------------------------------------------
// TAP Interface
//--------------------------------------------------
wire   [1:0]                    pad_sel_tap;
wire                            pad_tap_tck;
wire                            pad_tap_tms;
wire                            pad_tap_trst_n;
wire                            pad_tap_tdi;
wire                            pad_tap_tdo;

//--------------------------------------------------
// uC debugger TAP Interface
//--------------------------------------------------
wire                            pad_uc_tap_tck;
wire                            pad_uc_tap_tms;
wire                            pad_uc_tap_trst_n;
wire                            pad_uc_tap_tdi;
wire                            pad_uc_tap_tdo;

//--------------------------------------------------
// AUX/Sideband Interface
//--------------------------------------------------


//--------------------------------------------------
// PCS PIPE external Interface
//--------------------------------------------------
// *******************************
// Common pins
// *******************************
wire                            pad_pipe_clk_max;
wire                            pad_pipe_reset_n;
wire                            pad_pipe_rate;
wire                            pad_pipe_clk_max_req;
wire                            pad_pipe_clk_max_ack;
wire     [2-1:0]                pad_pipe_powerdown;
wire                            pad_pipe_pll0_en;
wire                            pad_pipe_pll0_ok;
wire                            pad_pma_cmn_ready;
wire                            pad_phy_interrupt;
wire                            pad_typec_conn_dir;
// *******************************
// Lane0 RX pins
// *******************************                        
wire                            pad_pipe_l00_rx_clk;
wire                            pad_pipe_l00_phy_status;
wire     [32-1:0]               pad_pipe_l00_rx_data;
wire     [8-1:0]                pad_pipe_l00_p2m_messagebus;
wire                            pad_pipe_l00_rx_start_block;
wire                            pad_pipe_l00_rx_data_valid;
wire                            pad_pipe_l00_rx_valid;
wire     [3-1:0]                pad_pipe_l00_rx_standby_status;
wire                            pad_pipe_l00_rx_elec_idle;
wire                            pad_pipe_l00_rx_standby;
wire                            pad_pipe_l00_rx_termination;
wire                            pad_pipe_l00_rx_eq_training;
// *******************************
// Lane0 TX pins
// *******************************              
wire                            pad_pipe_l00_clk;
wire     [32-1:0]               pad_pipe_l00_tx_data;
wire     [8-1:0]                pad_pipe_l00_m2p_messagebus;
wire                            pad_pipe_l00_tx_start_block;
wire                            pad_pipe_l00_tx_data_valid;
wire                            pad_pipe_l00_tx_det_rx_lpbk;
wire                            pad_pipe_l00_tx_elec_idle;
wire     [3-1:0]                pad_pipe_l00_powerdown;
wire     [2-1:0]                pad_pipe_l00_rate;
// *******************************
// Lane1 RX pins
// *******************************              
wire                            pad_pipe_l01_rx_clk;
wire                            pad_pipe_l01_phy_status;
wire     [32-1:0]               pad_pipe_l01_rx_data;
wire     [8-1:0]                pad_pipe_l01_p2m_messagebus;
wire                            pad_pipe_l01_rx_start_block;
wire                            pad_pipe_l01_rx_data_valid;
wire                            pad_pipe_l01_rx_valid;
wire     [3-1:0]                pad_pipe_l01_rx_standby_status;
wire                            pad_pipe_l01_rx_elec_idle;
wire                            pad_pipe_l01_rx_standby;
wire                            pad_pipe_l01_rx_termination;
wire                            pad_pipe_l01_rx_eq_training;
// *******************************
// Lane1 TX pins
// *******************************             
wire                            pad_pipe_l01_clk;
wire     [32-1:0]               pad_pipe_l01_tx_data;
wire     [8-1:0]                pad_pipe_l01_m2p_messagebus;
wire                            pad_pipe_l01_tx_start_block;
wire                            pad_pipe_l01_tx_data_valid;
wire                            pad_pipe_l01_tx_det_rx_lpbk;
wire                            pad_pipe_l01_tx_elec_idle;
wire     [3-1:0]                pad_pipe_l01_powerdown;
wire     [2-1:0]                pad_pipe_l01_rate;    

//----------------------------------------------------------------------
// Scan
//----------------------------------------------------------------------
wire          tie_scanmode   = 1'b0;
wire          tie_scanen     = 1'b0;
wire          tie_scanen_cg  = 1'b0;

/****************************************************************************\
|*                                                                          *|
|*      Functional Description                                              *|
|*                                                                          *|
\****************************************************************************/


//------------------------------------------------------------------------------
// MUX for Tap controllers
//------------------------------------------------------------------------------
tap_io_mux u_tap_io_mux (/*autoinst*/
        // Chip IO Interface
        .pad_sel_tap            (pad_sel_tap[1:0]               ), //input
        .pad_tap_tck            (pad_tap_tck                    ), //input
        .pad_tap_tms            (pad_tap_tms                    ), //input
        .pad_tap_trst_n         (pad_tap_trst_n                 ), //input
        .pad_tap_tdi            (pad_tap_tdi                    ), //input
        .pad_tap_tdo            (pad_tap_tdo                    ), //output
        // Shared
        .mux_tap_tck            (mux_tap_tck                    ), //output
        .mux_tap_trst_n         (mux_tap_trst_n                 ), //output
        .mux_tap_tdi            (mux_tap_tdi                    ), //output
        // TC JTAG
        .mux_tc_tap_tms         (mux_tc_tap_tms                 ), //output
        .mux_tc_tap_tdo         (mux_tc_tap_tdo                 ), //input
        // PHY JTAG
        .mux_tap_tms            (mux_tap_tms                    ), //output
        .mux_tap_tdo            (mux_tap_tdo                    )  //input
    );

testchip_tap2apb u_tap2apb(/*autoinst*/
        //Top level TAP pins
        .tap_tdi                (mux_tap_tdi                    ), //input
        .tap_tck                (mux_tap_tck                    ), //input
        .tap_tms                (mux_tc_tap_tms                 ), //input
        .tap_trst_n             (mux_tap_trst_n                 ), //input
        .tap_tdo                (mux_tc_tap_tdo                 ), //output
        .tap_tdoen              (/* unconnected */              ), //output
        // Top level NoC interface.
        .noc_clk                (pad_noc_clk                    ), //input
        .noc_reset_n            (pad_noc_reset_n                ), //input
        // CDB interface to NoC.
        .cdb_pclk               (cdb_pclk                       ), //output
        .cdb_preset_n           (cdb_preset_n                   ), //output
        .cdb_psel               (cdb_psel                       ), //output
        .cdb_penable            (cdb_penable                    ), //output
        .cdb_paddr              (cdb_paddr[31:0]                ), //output
        .cdb_pwrite             (cdb_pwrite                     ), //output
        .cdb_pwdata             (cdb_pwdata[31:0]               ), //output
        .cdb_prdata             (cdb_prdata[31:0]               ), //input
        .cdb_pready             (cdb_pready                     ), //input
        // Scan
        .scanmode               (tie_scanmode                   ), //input
        .scanen                 (tie_scanen                     ), //input
        .scanen_cg              (tie_scanen_cg                  )  //input
    );
//------------------------------------------------------------------------------
// TC clock and reset module
//------------------------------------------------------------------------------
testchip_clkrst u_tc_clkrst(/*autoinst*/
        //DDR clock
        .param_ddr_cal_cal_clk_div_sel      (param_ddr_cal_cal_clk_div_sel[3:0]         ), //input
        .param_ddr_pclk_div_sel             (param_ddr_pclk_div_sel[3:0]                ), //input
        .param_ddr_rx_pclk_en               (param_ddr_rx_pclk_en                       ), //input
        .ddr_cal_cal_clk                    (ddr_cal_cal_clk                            ), //output
        .ddr_pclk                           (ddr_pclk                                   ), //output
        .ddr_rx_pclk                        (ddr_rx_pclk                                ), //output
        // Scan
        .scanmode                           (tie_scanmode                               ), //input
        .scanen                             (tie_scanen                                 ), //input
        .scanen_cg                          (tie_scanen_cg                              ), //input
        //Clock
        .noc_clk                            (pad_noc_clk                                ), //input
        .uc_clk                             (pad_uc_clk                                 ), //input
        .cdb_pclk                           (cdb_pclk                                   ), //input
        .cmn_refclk0_int                    (pad_cmn_refclk0_int                        ), //input
        .cmn_refclk1_int                    (pad_cmn_refclk1_int                        ), //input
        //Reset
        .tc_reset_n                         (pad_tc_reset_n                             ), //input
        .noc_reset_n                        (pad_noc_reset_n                            ), //input
        .param_phy_ss_reset_n               (param_phy_ss_reset_n                       ), //input
        .param_pam3_ss_reset_n              (param_pam3_ss_reset_n                      ), //input
        .param_ddrio_ctrl_reset_n           (param_ddrio_ctrl_reset_n                   ), //input
        .param_test_clk_ctrl_reset_n        (param_test_clk_ctrl_reset_n                ), //input
        .phy_ss_reset_n                     (phy_ss_reset_n                             ), //output
        .pam3_ss_reset_n                    (pam3_ss_reset_n                            ), //output
        .ddrio_ctrl_reset_n                 (ddrio_ctrl_reset_n                         ), //output
        .test_clk_ctrl_reset_n              (test_clk_ctrl_reset_n                      ), //output
        .ddrio_ctrl_reset_n_sync            (ddrio_ctrl_reset_n_sync                    ), //output
        .ddr_pclk_reset_n_sync              (ddr_pclk_reset_n_sync                      ), //output
        // Test Clock
        .test_clk_phy                       (test_clk_phy                               ), //input
        .test_clk_pam3                      (test_clk_pam3                              ), //input
        .param_test_clk_sel                 (param_test_clk_sel[3:0]                    ), //input
        .param_test_clk_en                  (param_test_clk_en                          ), //input
        .test_clk                           (pad_test_clk                               ), //output
        //PHY Ref Clock
        `ifdef CDNS_PMA_PWR_AWARE 
        .avdd                               (avdd                                       ), //input
        .avdd_h                             (avdd_h                                     ), //input
        .gnd                                (gnd                                        ), //input
        `endif
        //TC REF CLK AUX 0
        //Analog Inputs	
        .tcauxda_0_ref_clk_p                (cmn_refclk0_p_phy                          ), //input
        .tcauxda_0_ref_clk_m                (cmn_refclk0_m_phy                          ), //input
        //Digital Inputs       
        .tcauxda_0_bg_start_hyst_dis        (param_tcauxda_0_bg_start_hyst_dis          ), //input
        .tcauxda_0_bg_start_adj             (param_tcauxda_0_bg_start_adj[1:0]          ), //input
        .tcauxda_0_bg_en                    (param_tcauxda_0_bg_en                      ), //input
        .tcauxda_0_bias_en                  (param_tcauxda_0_bias_en                    ), //input
        .tcauxda_0_bias_cur_adj             (param_tcauxda_0_bias_cur_adj[1:0]          ), //input
        .tcauxda_0_irext_trim               (param_tcauxda_0_irext_trim[5:0]            ), //input
        .tcauxda_0_pll_refclk_enable        (param_tcauxda_0_pll_refclk_enable          ), //input
        .tcauxda_0_ref_clk_int              (pad_cmn_refclk0_int                        ), //input
        .tcauxda_0_pll_refclk_sel           (param_tcauxda_0_pll_refclk_sel             ), //input
        .tcauxda_0_ref_clk0_ac_byp          (param_tcauxda_0_ref_clk0_ac_byp            ), //input
        .tcauxda_0_ref_clk0_dig_buf_en      (param_tcauxda_0_ref_clk0_dig_buf_en        ), //input
        .tcauxda_0_ref_clk0_dig_hyst_inc    (param_tcauxda_0_ref_clk0_dig_hyst_inc      ), //input
        .tcauxda_0_ref_clk0_filt_ctrl       (param_tcauxda_0_ref_clk0_filt_ctrl[1:0]    ), //input
        .tcauxda_0_ref_clk0_pll_buf_en      (param_tcauxda_0_ref_clk0_pll_buf_en        ), //input
        .tcauxda_0_ref_clk0_term_en         (param_tcauxda_0_ref_clk0_term_en           ), //input
        //Digital Outputs      
        .tcauxda_0_refclk_dig               (tcauxda_0_refclk_dig                       ), //output
        .tcauxda_0_pll_refclk_out           (tcauxda_0_pll_refclk_out                   ), //output
        //TC REF CLK AUX 1
        //Analog Inputs	
        .tcauxda_1_ref_clk_p                (cmn_refclk1_p_phy                          ), //input
        .tcauxda_1_ref_clk_m                (cmn_refclk1_m_phy                          ), //input
        //Digital Inputs       
        .tcauxda_1_bg_start_hyst_dis        (param_tcauxda_1_bg_start_hyst_dis          ), //input
        .tcauxda_1_bg_start_adj             (param_tcauxda_1_bg_start_adj[1:0]          ), //input
        .tcauxda_1_bg_en                    (param_tcauxda_1_bg_en                      ), //input
        .tcauxda_1_bias_en                  (param_tcauxda_1_bias_en                    ), //input
        .tcauxda_1_bias_cur_adj             (param_tcauxda_1_bias_cur_adj[1:0]          ), //input
        .tcauxda_1_irext_trim               (param_tcauxda_1_irext_trim[5:0]            ), //input
        .tcauxda_1_pll_refclk_enable        (param_tcauxda_1_pll_refclk_enable          ), //input
        .tcauxda_1_ref_clk_int              (pad_cmn_refclk1_int                        ), //input
        .tcauxda_1_pll_refclk_sel           (param_tcauxda_1_pll_refclk_sel             ), //input
        .tcauxda_1_ref_clk0_ac_byp          (param_tcauxda_1_ref_clk0_ac_byp            ), //input
        .tcauxda_1_ref_clk0_dig_buf_en      (param_tcauxda_1_ref_clk0_dig_buf_en        ), //input
        .tcauxda_1_ref_clk0_dig_hyst_inc    (param_tcauxda_1_ref_clk0_dig_hyst_inc      ), //input
        .tcauxda_1_ref_clk0_filt_ctrl       (param_tcauxda_1_ref_clk0_filt_ctrl[1:0]    ), //input
        .tcauxda_1_ref_clk0_pll_buf_en      (param_tcauxda_1_ref_clk0_pll_buf_en        ), //input
        .tcauxda_1_ref_clk0_term_en         (param_tcauxda_1_ref_clk0_term_en           ), //input
        //Digital Outputs      
        .tcauxda_1_refclk_dig               (tcauxda_1_refclk_dig                       ), //output
        .tcauxda_1_pll_refclk_out           (tcauxda_1_pll_refclk_out                   )  //output
    );

////------------------------------------------------------------------------------
//// TC registers module
////------------------------------------------------------------------------------
//testchip_top_reg_bank u_top_reg_bank(/*autoinst*/
//);
//

//------------------------------------------------------------------------------
// TC Noc Frabic
//------------------------------------------------------------------------------
usb4_tc_noc u_tc_noc(/*autoinst*/
        .tap2apb_pclk            (cdb_pclk                      ), //input
        .noc_clk                 (pad_noc_clk                   ), //input
        .rst_n                   (cdb_preset_n                  ), //input
        // apb_mstr
        .apb_mstr_paddr          (apb_mstr_paddr[31:0]          ), //input
        .apb_mstr_psel           (apb_mstr_psel                 ), //input
        .apb_mstr_penable        (apb_mstr_penable              ), //input
        .apb_mstr_pwrite         (apb_mstr_pwrite               ), //input
        .apb_mstr_pwdata         (apb_mstr_pwdata[31:0]         ), //input
        .apb_mstr_pstrb          (apb_mstr_pstrb[3:0]           ), //input
        .apb_mstr_pready         (apb_mstr_pready               ), //output
        .apb_mstr_prdata         (apb_mstr_prdata[31:0]         ), //output
        .apb_mstr_pslverr        (apb_mstr_pslverr              ), //output
        // cdb
        .cdb_paddr               (cdb_paddr[31:0]               ), //input
        .cdb_psel                (cdb_psel                      ), //input
        .cdb_penable             (cdb_penable                   ), //input
        .cdb_pwrite              (cdb_pwrite                    ), //input
        .cdb_pwdata              (cdb_pwdata[31:0]              ), //input
        .cdb_pstrb               (cdb_pstrb[3:0]                ), //input
        .cdb_pready              (cdb_pready                    ), //output
        .cdb_prdata              (cdb_prdata[31:0]              ), //output
        .cdb_pslverr             (cdb_pslverr                   ), //output
        // cmn_cdb
        .cmn_cdb_paddr           (cmn_cdb_paddr[8:0]            ), //output
        .cmn_cdb_psel            (cmn_cdb_psel                  ), //output
        .cmn_cdb_penable         (cmn_cdb_penable               ), //output
        .cmn_cdb_pwrite          (cmn_cdb_pwrite                ), //output
        .cmn_cdb_pwdata          (cmn_cdb_pwdata[31:0]          ), //output
        .cmn_cdb_pstrb           (cmn_cdb_pstrb[3:0]            ), //output
        .cmn_cdb_pready          (cmn_cdb_pready                ), //input
        .cmn_cdb_prdata          (cmn_cdb_prdata[31:0]          ), //input
        // tc_reg
        .tc_reg_paddr            (tc_reg_paddr[15:0]            ), //output
        .tc_reg_psel             (tc_reg_psel                   ), //output
        .tc_reg_penable          (tc_reg_penable                ), //output
        .tc_reg_pwrite           (tc_reg_pwrite                 ), //output
        .tc_reg_pwdata           (tc_reg_pwdata[31:0]           ), //output
        .tc_reg_pstrb            (tc_reg_pstrb[3:0]             ), //output
        .tc_reg_pready           (tc_reg_pready                 ), //input
        .tc_reg_prdata           (tc_reg_prdata[31:0]           ), //input
        // usb_sub_sys
        .usb_sub_sys_paddr       (usb_sub_sys_paddr[15:0]       ), //output
        .usb_sub_sys_psel        (usb_sub_sys_psel              ), //output
        .usb_sub_sys_penable     (usb_sub_sys_penable           ), //output
        .usb_sub_sys_pwrite      (usb_sub_sys_pwrite            ), //output
        .usb_sub_sys_pwdata      (usb_sub_sys_pwdata[31:0]      ), //output
        .usb_sub_sys_pstrb       (usb_sub_sys_pstrb[3:0]        ), //output
        .usb_sub_sys_pready      (usb_sub_sys_pready            ), //input
        .usb_sub_sys_prdata      (usb_sub_sys_prdata[31:0]      ), //input
        // pam3_sub_sys
        .pam3_sub_sys_paddr      (pam3_sub_sys_paddr[15:0]      ), //output
        .pam3_sub_sys_psel       (pam3_sub_sys_psel             ), //output
        .pam3_sub_sys_penable    (pam3_sub_sys_penable          ), //output
        .pam3_sub_sys_pwrite     (pam3_sub_sys_pwrite           ), //output
        .pam3_sub_sys_pwdata     (pam3_sub_sys_pwdata[31:0]     ), //output
        .pam3_sub_sys_pstrb      (pam3_sub_sys_pstrb[3:0]       ), //output
        .pam3_sub_sys_pready     (pam3_sub_sys_pready           ), //input
        .pam3_sub_sys_prdata     (pam3_sub_sys_prdata[31:0]     ), //input
        // apb_tgt
        .apb_tgt_paddr           (apb_tgt_paddr[17:0]           ), //output
        .apb_tgt_psel            (apb_tgt_psel                  ), //output
        .apb_tgt_penable         (apb_tgt_penable               ), //output
        .apb_tgt_pwrite          (apb_tgt_pwrite                ), //output
        .apb_tgt_pwdata          (apb_tgt_pwdata[31:0]          ), //output
        .apb_tgt_pstrb           (apb_tgt_pstrb[3:0]            ), //output
        .apb_tgt_pready          (apb_tgt_pready                ), //input
        .apb_tgt_prdata          (apb_tgt_prdata[31:0]          ), //input
        .apb_tgt_pslverr         (apb_tgt_pslverr               ), //input
        // xcvr_ln_0
        .xcvr_ln_0_paddr         (xcvr_ln_0_paddr[9:0]          ), //output
        .xcvr_ln_0_psel          (xcvr_ln_0_psel                ), //output
        .xcvr_ln_0_penable       (xcvr_ln_0_penable             ), //output
        .xcvr_ln_0_pwrite        (xcvr_ln_0_pwrite              ), //output
        .xcvr_ln_0_pwdata        (xcvr_ln_0_pwdata[31:0]        ), //output
        .xcvr_ln_0_pstrb         (xcvr_ln_0_pstrb[3:0]          ), //output
        .xcvr_ln_0_pready        (xcvr_ln_0_pready              ), //input
        .xcvr_ln_0_prdata        (xcvr_ln_0_prdata[31:0]        )  //input
    );

//------------------------------------------------------------------------------
// MUX for UC Denug Tap controllers
//------------------------------------------------------------------------------
tap_io_mux_dbgr u_tap_io_mux_dbgr(/*autoinst*/
        // Chip IO Interface
        .param_uc_sel_tap       (param_uc_sel_tap[3:0]          ), //input
        .pad_uc_tap_tck         (pad_uc_tap_tck                 ), //input
        .pad_uc_tap_tms         (pad_uc_tap_tms                 ), //input
        .pad_uc_tap_trst_n      (pad_uc_tap_trst_n              ), //input
        .pad_uc_tap_tdi         (pad_uc_tap_tdi                 ), //input
        .pad_uc_tap_tdo         (pad_uc_tap_tdo                 ), //output
        // uC debugger JTAG interfaces for x1 and x2 PHY 
        // Shared signals
        .mux_uc_tap_tck         (mux_uc_tap_tck                 ), //output
        .mux_uc_tap_trst        (mux_uc_tap_trst                ), //output
        .mux_uc_tap_tdi         (mux_uc_tap_tdi                 ), //output
        // x2 PHY lane 0 uC
        .mux_uc_l01_tap_tms     (mux_uc_l01_tap_tms             ), //output
        .mux_uc_l01_tap_tdo     (mux_uc_l01_tap_tdo             ), //input
        // x2 PHY lane 1 uC
        .mux_uc_l23_tap_tms     (mux_uc_l23_tap_tms             ), //output
        .mux_uc_l23_tap_tdo     (mux_uc_l23_tap_tdo             ), //input
        // x2 PHY top uC
        .mux_uc_top_tap_tms     (mux_uc_top_tap_tms             ), //output
        .mux_uc_top_tap_tdo     (mux_uc_top_tap_tdo             )  //input
    );

//------------------------------------------------------------------------------
// USB Type-C PHY sub-system
//------------------------------------------------------------------------------
phy_subsystem u_phy_subsystem(/*autoinst*/
        //--------------------------------------------------
        // Supply/Ground Pads
        //--------------------------------------------------
        `ifdef CDNS_PHY_PWR_AWARE // @RELEASE@
        // *******************************
        // PHY Power pins
        // *******************************
        .agnd                          (agnd                                     ), //input
        .avdd_clk                      (avdd_clk                                 ), //input
        .avdd_h                        (avdd_h                                   ), //input
        .avdd                          (avdd                                     ), //input
        .avdd_tx0                      (avdd_tx0                                 ), //input
        .avdd_tx1                      (avdd_tx1                                 ), //input
        .avdd_tx2                      (avdd_tx2                                 ), //input
        .avdd_tx3                      (avdd_tx3                                 ), //input
        .avdd_rx                       (avdd_rx                                  ), //input
        .cmn_aonvdd                    (cmn_aonvdd                               ), //input
        .vdd                           (vdd                                      ), //input
        `endif // @RELEASE@
        // Scan
        .scanmode                      (tie_scanmode                             ), //input
        .scanen                        (tie_scanen                               ), //input
        .scanen_cg                     (tie_scanen_cg                            ), //input
        //--------------------------------------------------
        // System Clocks
        //--------------------------------------------------
        .cmn_refclk0_int               (tcauxda_0_pll_refclk_out                 ), //input
        .cmn_refclk1_int               (tcauxda_1_pll_refclk_out                 ), //input
        //--------------------------------------------------
        // uC clock
        //--------------------------------------------------
        .uc_clk                        (pad_uc_clk                               ), //input
        //--------------------------------------------------
        // Sub-system reset
        //--------------------------------------------------
        .reset_n                       (phy_ss_reset_n                           ), //input
        //--------------------------------------------------
        // PMA External Interface
        // MP PHY Interface
        //--------------------------------------------------
        .xcvr_p_ln_0                   (xcvr_p_ln_0_phy                          ), //inout
        .xcvr_m_ln_0                   (xcvr_m_ln_0_phy                          ), //inout
        .xcvr_p_ln_1                   (xcvr_p_ln_1_phy                          ), //inout
        .xcvr_m_ln_1                   (xcvr_m_ln_1_phy                          ), //inout
        .xcvr_p_ln_2                   (xcvr_p_ln_2_phy                          ), //inout
        .xcvr_m_ln_2                   (xcvr_m_ln_2_phy                          ), //inout
        .xcvr_p_ln_3                   (xcvr_p_ln_3_phy                          ), //inout
        .xcvr_m_ln_3                   (xcvr_m_ln_3_phy                          ), //inout
        .cmn_rext                      (cmn_rext_phy                             ), //input
        //--------------------------------------------------
        //Test Interface
        //--------------------------------------------------
        .atb_0                         (atb_0_phy                                ), //inout
        .atb_1                         (atb_1_phy                                ), //inout
        .param_dtb_data_sel            (param_dtb_data_sel[3:0]                  ), //input
        .param_dtb_data_en             (param_dtb_data_en                        ), //input
        .dtb_data_pam3                 (dtb_data_pam3[31:0]                      ), //input
        .dtb_data_tc                   (dtb_data_tc[31:0]                        ), //input
        .test_clk                      (test_clk_phy                             ), //output
        //--------------------------------------------------
        // TAP Interface
        //--------------------------------------------------
        .tap_tck                       (mux_tap_tck                              ), //input
        .tap_tms                       (mux_tap_tms                              ), //input
        .tap_trst_n                    (mux_tap_trst_n                           ), //input
        .tap_tdi                       (mux_tap_tdi                              ), //input
        .tap_tdo                       (mux_tap_tdo                              ), //output
        .tap_tdoen                     (/* unconnected */                        ), //output
        //--------------------------------------------------
        // uC debugger TAP Interface
        //--------------------------------------------------
        `ifdef CDN_TESTCHIP_UC_DBGR
        //uC debugger Tap interfaces
        .uc_top_tap_tck                (mux_uc_tap_tck                           ), //input
        .uc_top_tap_tms                (mux_uc_top_tap_tms                       ), //input
        .uc_top_tap_trst_n             (mux_uc_tap_trst_n                        ), //input
        .uc_top_tap_tdi                (mux_uc_tap_tdi                           ), //input
        .uc_top_tap_tdo                (mux_uc_top_tap_tdo                       ), //output
        .uc_top_tap_tdoen              (/* unconnected */                        ), //output
        `ifndef CDN_MPPHY_LANE_UC_RMV
        .uc_l01_tap_tck                (mux_uc_tap_tck                           ), //input
        .uc_l01_tap_tms                (mux_uc_l01_tap_tms                       ), //input
        .uc_l01_tap_trst_n             (mux_uc_tap_trst_n                        ), //input
        .uc_l01_tap_tdi                (mux_uc_tap_tdi                           ), //input
        .uc_l01_tap_tdo                (mux_uc_l01_tap_tdo                       ), //output
        .uc_l01_tap_tdoen              (/* unconnected */                        ), //output
        .uc_l23_tap_tck                (mux_uc_tap_tck                           ), //input
        .uc_l23_tap_tms                (mux_uc_l23_tap_tms                       ), //input
        .uc_l23_tap_trst_n             (mux_uc_tap_trst_n                        ), //input
        .uc_l23_tap_tdi                (mux_uc_tap_tdi                           ), //input
        .uc_l23_tap_tdo                (mux_uc_l23_tap_tdo                       ), //output
        .uc_l23_tap_tdoen              (/* unconnected */                        ), //output
        `endif
        `endif
        //--------------------------------------------------
        // APB Interface
        //--------------------------------------------------
        // *******************************
        // External APB target interface
        // *******************************
        .apb_pclk                      (pad_noc_clk                              ), //input
        .apb_preset_n                  (cdb_preset_n                             ), //input
        .apb_tgt_penable               (apb_tgt_penable                          ), //input
        .apb_tgt_psel                  (apb_tgt_psel                             ), //input
        .apb_tgt_pwrite                (apb_tgt_pwrite                           ), //input
        .apb_tgt_paddr                 (apb_tgt_paddr[17:0]                      ), //input
        .apb_tgt_pwdata                (apb_tgt_pwdata[31:0]                     ), //input
        .apb_tgt_prdata                (apb_tgt_prdata[31:0]                     ), //output
        .apb_tgt_pready                (apb_tgt_pready                           ), //output
        .apb_tgt_perr                  (apb_tgt_pslverr                          ), //output
        // *******************************
        // External APB master interface
        // *******************************
        .apb_mstr_penable              (apb_mstr_penable                         ), //output
        .apb_mstr_psel                 (apb_mstr_psel                            ), //output
        .apb_mstr_pwrite               (apb_mstr_pwrite                          ), //output
        .apb_mstr_paddr                (apb_mstr_paddr[31:0]                     ), //output
        .apb_mstr_pwdata               (apb_mstr_pwdata[31:0]                    ), //output
        .apb_mstr_prdata               (apb_mstr_prdata[31:0]                    ), //input
        .apb_mstr_pready               (apb_mstr_pready                          ), //input
        .apb_mstr_perr                 (apb_mstr_pslverr                         ), //input
        // *******************************
        // Subsystem APB master interface
        // *******************************
        .usb_sub_sys_pclk              (pad_noc_clk                              ), //input
        .usb_sub_sys_preset_n          (cdb_preset_n                             ), //input
        .usb_sub_sys_penable           (usb_sub_sys_penable                      ), //input
        .usb_sub_sys_psel              (usb_sub_sys_psel                         ), //input
        .usb_sub_sys_pwrite            (usb_sub_sys_pwrite                       ), //input
        .usb_sub_sys_paddr             (usb_sub_sys_paddr[15:0]                  ), //input
        .usb_sub_sys_pwdata            (usb_sub_sys_pwdata[31:0]                 ), //input
        .usb_sub_sys_prdata            (usb_sub_sys_prdata[31:0]                 ), //output
        .usb_sub_sys_pready            (usb_sub_sys_pready                       ), //output
        //--------------------------------------------------
        // PCS PIPE external Interface
        //--------------------------------------------------
        // *******************************
        // Common pins
        // *******************************
        .pipe_clk_max                  (pad_pipe_clk_max                         ), //output
        .pipe_reset_n                  (pad_pipe_reset_n                         ), //input
        .pipe_rate                     (pad_pipe_rate                            ), //input
        .pipe_clk_max_req              (pad_pipe_clk_max_req                     ), //input
        .pipe_clk_max_ack              (pad_pipe_clk_max_ack                     ), //output
        .pipe_powerdown                (pad_pipe_powerdown[2-1:0]                ), //input
        .pipe_pll0_en                  (pad_pipe_pll0_en                         ), //input
        .pipe_pll0_ok                  (pad_pipe_pll0_ok                         ), //output
        .pma_cmn_ready                 (pad_pma_cmn_ready                        ), //output
        .phy_interrupt                 (pad_phy_interrupt                        ), //output
        .typec_conn_dir                (pad_typec_conn_dir                       ), //input
        // *******************************
        // Lane0 RX pins
        // *******************************                        
        .pipe_l00_rx_clk               (pad_pipe_l00_rx_clk                      ), //output
        .pipe_l00_phy_status           (pad_pipe_l00_phy_status                  ), //output
        .pipe_l00_rx_data              (pad_pipe_l00_rx_data[32-1:0]             ), //output
        .pma_tx_td_ln_0                (pad_pma_tx_td_ln_0[32-1:0]               ), //input
        .pipe_l00_p2m_messagebus       (pad_pipe_l00_p2m_messagebus[8-1:0]       ), //output
        .pipe_l00_rx_start_block       (pad_pipe_l00_rx_start_block              ), //output
        .pipe_l00_rx_data_valid        (pad_pipe_l00_rx_data_valid               ), //output
        .pma_tx_elec_idle_ln_0         (pad_pma_tx_elec_idle_ln_0                ), //input
        .pipe_l00_rx_valid             (pad_pipe_l00_rx_valid                    ), //output
        .pipe_l00_rx_standby_status    (pad_pipe_l00_rx_standby_status[3-1:0]    ), //output
        .pipe_l00_rx_elec_idle         (pad_pipe_l00_rx_elec_idle                ), //output
        .pipe_l00_rx_standby           (pad_pipe_l00_rx_standby                  ), //input
        .pipe_l00_rx_termination       (pad_pipe_l00_rx_termination              ), //input
        .pipe_l00_rx_eq_training       (pad_pipe_l00_rx_eq_training              ), //input
        // *******************************
        // Lane0 TX pins
        // *******************************              
        .pipe_l00_clk                  (pad_pipe_l00_clk                         ), //input
        .pipe_l00_tx_data              (pad_pipe_l00_tx_data[32-1:0]             ), //input
        .pipe_l00_m2p_messagebus       (pad_pipe_l00_m2p_messagebus[8-1:0]       ), //input
        .pipe_l00_tx_start_block       (pad_pipe_l00_tx_start_block              ), //input
        .pipe_l00_tx_data_valid        (pad_pipe_l00_tx_data_valid               ), //input
        .pipe_l00_tx_det_rx_lpbk       (pad_pipe_l00_tx_det_rx_lpbk              ), //input
        .pipe_l00_tx_elec_idle         (pad_pipe_l00_tx_elec_idle                ), //input
        .pipe_l00_powerdown            (pad_pipe_l00_powerdown[3-1:0]            ), //input
        .pipe_l00_rate                 (pad_pipe_l00_rate[2-1:0]                 ), //input
        // *******************************
        // Lane1 RX pins
        // *******************************              
        .pipe_l01_rx_clk               (pad_pipe_l01_rx_clk                      ), //output
        .pipe_l01_phy_status           (pad_pipe_l01_phy_status                  ), //output
        .pipe_l01_rx_data              (pad_pipe_l01_rx_data[32-1:0]             ), //output
        .pma_tx_td_ln_1                (pad_pma_tx_td_ln_1[32-1:0]               ), //input
        .pipe_l01_p2m_messagebus       (pad_pipe_l01_p2m_messagebus[8-1:0]       ), //output
        .pipe_l01_rx_start_block       (pad_pipe_l01_rx_start_block              ), //output
        .pipe_l01_rx_data_valid        (pad_pipe_l01_rx_data_valid               ), //output
        .pma_tx_elec_idle_ln_0         (pad_pma_tx_elec_idle_ln_0                ), //input
        .pipe_l01_rx_valid             (pad_pipe_l01_rx_valid                    ), //output
        .pipe_l01_rx_standby_status    (pad_pipe_l01_rx_standby_status[3-1:0]    ), //output
        .pipe_l01_rx_elec_idle         (pad_pipe_l01_rx_elec_idle                ), //output
        .pipe_l01_rx_standby           (pad_pipe_l01_rx_standby                  ), //input
        .pipe_l01_rx_termination       (pad_pipe_l01_rx_termination              ), //input
        .pipe_l01_rx_eq_training       (pad_pipe_l01_rx_eq_training              ), //input
        // *******************************
        // Lane1 TX pins
        // *******************************             
        .pipe_l01_clk                  (pad_pipe_l01_clk                         ), //input
        .pipe_l01_tx_data              (pad_pipe_l01_tx_data[32-1:0]             ), //input
        .pipe_l01_m2p_messagebus       (pad_pipe_l01_m2p_messagebus[8-1:0]       ), //input
        .pipe_l01_tx_start_block       (pad_pipe_l01_tx_start_block              ), //input
        .pipe_l01_tx_data_valid        (pad_pipe_l01_tx_data_valid               ), //input
        .pipe_l01_tx_det_rx_lpbk       (pad_pipe_l01_tx_det_rx_lpbk              ), //input
        .pipe_l01_tx_elec_idle         (pad_pipe_l01_tx_elec_idle                ), //input
        .pipe_l01_powerdown            (pad_pipe_l01_powerdown[3-1:0]            ), //input
        .pipe_l01_rate                 (pad_pipe_l01_rate[2-1:0]                 )  //input
    );

//------------------------------------------------------------------------------
// PAM3 PMA sub-system
//------------------------------------------------------------------------------
pam3_subsystem u_pam3_subsystem(/*autoinst*/
        // Top level bump signals.
        `ifdef CDNS_PMA_PWR_AWARE // @RELEASE@
        .agnd                     (agnd                         ), //input
        .avdd_clk                 (avdd_clk                     ), //input
        .avdd_h                   (avdd_h                       ), //input
        .avdd                     (avdd                         ), //input
        .avdd_tx0                 (avdd_tx0                     ), //input
        .avdd_tx1                 (avdd_tx1                     ), //input
        .avdd_tx2                 (avdd_tx2                     ), //input
        .avdd_tx3                 (avdd_tx3                     ), //input
        .avdd_rx                  (avdd_rx                      ), //input
        .cmn_aonvdd               (cmn_aonvdd                   ), //input
        .vdd                      (vdd                          ), //input
        `endif // @RELEASE@
        // Scan
        .scanmode                 (tie_scanmode                 ), //input
        .scanen                   (tie_scanen                   ), //input
        .scanen_cg                (tie_scanen_cg                ), //input
        //Clock   
        .cmn_ref_clk0_int         (pad_cmn_refclk0_int          ), //input
        .cmn_ref_clk1_int         (pad_cmn_refclk1_int          ), //input
        .cmn_refclk0_p            (cmn_refclk0_p_pam3           ), //input
        .cmn_refclk0_m            (cmn_refclk0_m_pam3           ), //input
        .cmn_refclk1_p            (cmn_refclk1_p_pam3           ), //input
        .cmn_refclk1_m            (cmn_refclk1_m_pam3           ), //input
        // Sub-system reset
        .reset_n                  (pam3_ss_reset_n              ), //input
        // PMA common CDB signals.
        .cmn_cdb_pclk             (pad_noc_clk                  ), //input
        .cmn_cdb_preset_n         (cdb_preset_n                 ), //input
        .cmn_cdb_penable          (cmn_cdb_penable              ), //input
        .cmn_cdb_psel             (cmn_cdb_psel                 ), //input
        .cmn_cdb_paddr            (cmn_cdb_paddr[8:0]           ), //input
        .cmn_cdb_pwrite           (cmn_cdb_pwrite               ), //input
        .cmn_cdb_pwdata           (cmn_cdb_pwdata[31:0]         ), //input
        .cmn_cdb_prdata           (cmn_cdb_prdata[31:0]         ), //output
        .cmn_cdb_pready           (cmn_cdb_pready               ), //output
        // PMA Transceiver CDB signals.
        .xcvr_ln_0_pclk           (pad_noc_clk                  ), //input
        .xcvr_ln_0_preset_n       (cdb_preset_n                 ), //input
        .xcvr_ln_0_penable        (xcvr_ln_0_penable            ), //input
        .xcvr_ln_0_psel           (xcvr_ln_0_psel               ), //input
        .xcvr_ln_0_paddr          (xcvr_ln_0_paddr[9:0]         ), //input
        .xcvr_ln_0_pwrite         (xcvr_ln_0_pwrite             ), //input
        .xcvr_ln_0_pwdata         (xcvr_ln_0_pwdata[31:0]       ), //input
        .xcvr_ln_0_prdata         (xcvr_ln_0_prdata[31:0]       ), //output
        .xcvr_ln_0_pready         (xcvr_ln_0_pready             ), //output
        // PAM3 sub system CDB signals.
        .pam3_sub_sys_pclk        (pad_noc_clk                  ), //input
        .pam3_sub_sys_preset_n    (cdb_preset_n                 ), //input
        .pam3_sub_sys_paddr       (pam3_sub_sys_paddr[15:0]     ), //input
        .pam3_sub_sys_psel        (pam3_sub_sys_psel            ), //input
        .pam3_sub_sys_penable     (pam3_sub_sys_penable         ), //input
        .pam3_sub_sys_pwrite      (pam3_sub_sys_pwrite          ), //input
        .pam3_sub_sys_pwdata      (pam3_sub_sys_pwdata[31:0]    ), //input
        .pam3_sub_sys_pstrb       (pam3_sub_sys_pstrb[3:0]      ), //input
        .pam3_sub_sys_pready      (pam3_sub_sys_pready          ), //output
        .pam3_sub_sys_prdata      (pam3_sub_sys_prdata[31:0]    ), //output
        //BUMP
        .cmn_rext                 (cmn_rext_pam3                ), //inout
        .xcvr_p_ln_0              (xcvr_p_ln_0_pam3             ), //inout
        .xcvr_m_ln_0              (xcvr_m_ln_0_pam3             ), //inout
        // Digital Test Bus   
        `ifndef CDN_MPPHY_RMV_DTB // @RELEASE@
        .dtb_data                 (dtb_data_pam3[31:0]          ), //output
        .dtb_clk                  (dtb_clk_pam3                 ), //output
        `endif // @RELEASE@   
        //ATB
        .cmn_atb_core_0           (atb_0_pam3                   ), //inout
        .cmn_atb_core_1           (atb_1_pam3                   )  //inout
    );

////------------------------------------------------------------------------------
//// Test Chip Pads
////------------------------------------------------------------------------------
//module testchip_pads (/*autoinst*/
//);


endmodule

// Local Variables:
// verilog-library-directories:(".")
// verilog-library-directories:("./phy_subsystem")
// verilog-library-directories:("./pam3_subsystem")
// verilog-library-directories:("./noc/usb4_tc_noc/rtl/noc")
// End:

