`include"cdn_message_bus_sequence.sv"
