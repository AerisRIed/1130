`include"cdn_alt_mode_phy_test_base.sv"


