`include "cdn_phy_bring_up_test_base.sv"