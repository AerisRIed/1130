`include"cdn_u4_pcie_base_sequence.sv"


