`ifndef GATESIM__SV
`define GATESIM__SV
//TODO gatesim issue like:
    //initial value of memory

    //sdf anno

    //other tie_offs

    //no timing check

    //other block needed

`endif