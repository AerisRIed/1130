interface cdn_jtag_1687_interface(input tck);

logic tdo;
logic trst = 0;
logic clockdr;
logic shiftdr;
logic updatedr;
logic capturedr;
logic instruction_decode_instr_1;
logic instruction_decode_instr_2;
logic instruction_decode_instr_3;
logic instruction_decode_instr_4;
logic instruction_decode_instr_5;
endinterface
