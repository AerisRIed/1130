`include"cdn_u4_vip_base_sequence.sv"
